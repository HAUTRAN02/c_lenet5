// tb.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module tb (
	);

	wire  [63:0] avgpooling1_inst_avmm_0_rw_readdata;                                                           // mm_agent_dpi_bfm_avgpooling1_avmm_0_rw_inst:avs_readdata -> avgpooling1_inst:avmm_0_rw_readdata
	wire  [63:0] avgpooling1_inst_avmm_0_rw_address;                                                            // avgpooling1_inst:avmm_0_rw_address -> mm_agent_dpi_bfm_avgpooling1_avmm_0_rw_inst:avs_address
	wire   [7:0] avgpooling1_inst_avmm_0_rw_byteenable;                                                         // avgpooling1_inst:avmm_0_rw_byteenable -> mm_agent_dpi_bfm_avgpooling1_avmm_0_rw_inst:avs_byteenable
	wire         avgpooling1_inst_avmm_0_rw_read;                                                               // avgpooling1_inst:avmm_0_rw_read -> mm_agent_dpi_bfm_avgpooling1_avmm_0_rw_inst:avs_read
	wire         avgpooling1_inst_avmm_0_rw_write;                                                              // avgpooling1_inst:avmm_0_rw_write -> mm_agent_dpi_bfm_avgpooling1_avmm_0_rw_inst:avs_write
	wire  [63:0] avgpooling1_inst_avmm_0_rw_writedata;                                                          // avgpooling1_inst:avmm_0_rw_writedata -> mm_agent_dpi_bfm_avgpooling1_avmm_0_rw_inst:avs_writedata
	wire  [63:0] avgpooling2_inst_avmm_0_rw_readdata;                                                           // mm_agent_dpi_bfm_avgpooling2_avmm_0_rw_inst:avs_readdata -> avgpooling2_inst:avmm_0_rw_readdata
	wire  [63:0] avgpooling2_inst_avmm_0_rw_address;                                                            // avgpooling2_inst:avmm_0_rw_address -> mm_agent_dpi_bfm_avgpooling2_avmm_0_rw_inst:avs_address
	wire   [7:0] avgpooling2_inst_avmm_0_rw_byteenable;                                                         // avgpooling2_inst:avmm_0_rw_byteenable -> mm_agent_dpi_bfm_avgpooling2_avmm_0_rw_inst:avs_byteenable
	wire         avgpooling2_inst_avmm_0_rw_read;                                                               // avgpooling2_inst:avmm_0_rw_read -> mm_agent_dpi_bfm_avgpooling2_avmm_0_rw_inst:avs_read
	wire         avgpooling2_inst_avmm_0_rw_write;                                                              // avgpooling2_inst:avmm_0_rw_write -> mm_agent_dpi_bfm_avgpooling2_avmm_0_rw_inst:avs_write
	wire  [63:0] avgpooling2_inst_avmm_0_rw_writedata;                                                          // avgpooling2_inst:avmm_0_rw_writedata -> mm_agent_dpi_bfm_avgpooling2_avmm_0_rw_inst:avs_writedata
	wire  [63:0] conv1_inst_avmm_0_rw_readdata;                                                                 // mm_agent_dpi_bfm_conv1_avmm_0_rw_inst:avs_readdata -> conv1_inst:avmm_0_rw_readdata
	wire  [63:0] conv1_inst_avmm_0_rw_address;                                                                  // conv1_inst:avmm_0_rw_address -> mm_agent_dpi_bfm_conv1_avmm_0_rw_inst:avs_address
	wire   [7:0] conv1_inst_avmm_0_rw_byteenable;                                                               // conv1_inst:avmm_0_rw_byteenable -> mm_agent_dpi_bfm_conv1_avmm_0_rw_inst:avs_byteenable
	wire         conv1_inst_avmm_0_rw_read;                                                                     // conv1_inst:avmm_0_rw_read -> mm_agent_dpi_bfm_conv1_avmm_0_rw_inst:avs_read
	wire         conv1_inst_avmm_0_rw_write;                                                                    // conv1_inst:avmm_0_rw_write -> mm_agent_dpi_bfm_conv1_avmm_0_rw_inst:avs_write
	wire  [63:0] conv1_inst_avmm_0_rw_writedata;                                                                // conv1_inst:avmm_0_rw_writedata -> mm_agent_dpi_bfm_conv1_avmm_0_rw_inst:avs_writedata
	wire  [63:0] conv2_inst_avmm_0_rw_readdata;                                                                 // mm_agent_dpi_bfm_conv2_avmm_0_rw_inst:avs_readdata -> conv2_inst:avmm_0_rw_readdata
	wire  [63:0] conv2_inst_avmm_0_rw_address;                                                                  // conv2_inst:avmm_0_rw_address -> mm_agent_dpi_bfm_conv2_avmm_0_rw_inst:avs_address
	wire   [7:0] conv2_inst_avmm_0_rw_byteenable;                                                               // conv2_inst:avmm_0_rw_byteenable -> mm_agent_dpi_bfm_conv2_avmm_0_rw_inst:avs_byteenable
	wire         conv2_inst_avmm_0_rw_read;                                                                     // conv2_inst:avmm_0_rw_read -> mm_agent_dpi_bfm_conv2_avmm_0_rw_inst:avs_read
	wire         conv2_inst_avmm_0_rw_write;                                                                    // conv2_inst:avmm_0_rw_write -> mm_agent_dpi_bfm_conv2_avmm_0_rw_inst:avs_write
	wire  [63:0] conv2_inst_avmm_0_rw_writedata;                                                                // conv2_inst:avmm_0_rw_writedata -> mm_agent_dpi_bfm_conv2_avmm_0_rw_inst:avs_writedata
	wire  [63:0] fc1_inst_avmm_0_rw_readdata;                                                                   // mm_agent_dpi_bfm_fc1_avmm_0_rw_inst:avs_readdata -> fc1_inst:avmm_0_rw_readdata
	wire  [63:0] fc1_inst_avmm_0_rw_address;                                                                    // fc1_inst:avmm_0_rw_address -> mm_agent_dpi_bfm_fc1_avmm_0_rw_inst:avs_address
	wire   [7:0] fc1_inst_avmm_0_rw_byteenable;                                                                 // fc1_inst:avmm_0_rw_byteenable -> mm_agent_dpi_bfm_fc1_avmm_0_rw_inst:avs_byteenable
	wire         fc1_inst_avmm_0_rw_read;                                                                       // fc1_inst:avmm_0_rw_read -> mm_agent_dpi_bfm_fc1_avmm_0_rw_inst:avs_read
	wire         fc1_inst_avmm_0_rw_write;                                                                      // fc1_inst:avmm_0_rw_write -> mm_agent_dpi_bfm_fc1_avmm_0_rw_inst:avs_write
	wire  [63:0] fc1_inst_avmm_0_rw_writedata;                                                                  // fc1_inst:avmm_0_rw_writedata -> mm_agent_dpi_bfm_fc1_avmm_0_rw_inst:avs_writedata
	wire  [63:0] fc3_inst_avmm_0_rw_readdata;                                                                   // mm_agent_dpi_bfm_fc3_avmm_0_rw_inst:avs_readdata -> fc3_inst:avmm_0_rw_readdata
	wire  [63:0] fc3_inst_avmm_0_rw_address;                                                                    // fc3_inst:avmm_0_rw_address -> mm_agent_dpi_bfm_fc3_avmm_0_rw_inst:avs_address
	wire   [7:0] fc3_inst_avmm_0_rw_byteenable;                                                                 // fc3_inst:avmm_0_rw_byteenable -> mm_agent_dpi_bfm_fc3_avmm_0_rw_inst:avs_byteenable
	wire         fc3_inst_avmm_0_rw_read;                                                                       // fc3_inst:avmm_0_rw_read -> mm_agent_dpi_bfm_fc3_avmm_0_rw_inst:avs_read
	wire         fc3_inst_avmm_0_rw_write;                                                                      // fc3_inst:avmm_0_rw_write -> mm_agent_dpi_bfm_fc3_avmm_0_rw_inst:avs_write
	wire  [63:0] fc3_inst_avmm_0_rw_writedata;                                                                  // fc3_inst:avmm_0_rw_writedata -> mm_agent_dpi_bfm_fc3_avmm_0_rw_inst:avs_writedata
	wire  [63:0] relu1_inst_avmm_0_rw_readdata;                                                                 // mm_agent_dpi_bfm_relu1_avmm_0_rw_inst:avs_readdata -> relu1_inst:avmm_0_rw_readdata
	wire  [63:0] relu1_inst_avmm_0_rw_address;                                                                  // relu1_inst:avmm_0_rw_address -> mm_agent_dpi_bfm_relu1_avmm_0_rw_inst:avs_address
	wire   [7:0] relu1_inst_avmm_0_rw_byteenable;                                                               // relu1_inst:avmm_0_rw_byteenable -> mm_agent_dpi_bfm_relu1_avmm_0_rw_inst:avs_byteenable
	wire         relu1_inst_avmm_0_rw_read;                                                                     // relu1_inst:avmm_0_rw_read -> mm_agent_dpi_bfm_relu1_avmm_0_rw_inst:avs_read
	wire         relu1_inst_avmm_0_rw_write;                                                                    // relu1_inst:avmm_0_rw_write -> mm_agent_dpi_bfm_relu1_avmm_0_rw_inst:avs_write
	wire  [63:0] relu1_inst_avmm_0_rw_writedata;                                                                // relu1_inst:avmm_0_rw_writedata -> mm_agent_dpi_bfm_relu1_avmm_0_rw_inst:avs_writedata
	wire  [63:0] relu2_inst_avmm_0_rw_readdata;                                                                 // mm_agent_dpi_bfm_relu2_avmm_0_rw_inst:avs_readdata -> relu2_inst:avmm_0_rw_readdata
	wire  [63:0] relu2_inst_avmm_0_rw_address;                                                                  // relu2_inst:avmm_0_rw_address -> mm_agent_dpi_bfm_relu2_avmm_0_rw_inst:avs_address
	wire   [7:0] relu2_inst_avmm_0_rw_byteenable;                                                               // relu2_inst:avmm_0_rw_byteenable -> mm_agent_dpi_bfm_relu2_avmm_0_rw_inst:avs_byteenable
	wire         relu2_inst_avmm_0_rw_read;                                                                     // relu2_inst:avmm_0_rw_read -> mm_agent_dpi_bfm_relu2_avmm_0_rw_inst:avs_read
	wire         relu2_inst_avmm_0_rw_write;                                                                    // relu2_inst:avmm_0_rw_write -> mm_agent_dpi_bfm_relu2_avmm_0_rw_inst:avs_write
	wire  [63:0] relu2_inst_avmm_0_rw_writedata;                                                                // relu2_inst:avmm_0_rw_writedata -> mm_agent_dpi_bfm_relu2_avmm_0_rw_inst:avs_writedata
	wire  [63:0] relu3_inst_avmm_0_rw_readdata;                                                                 // mm_agent_dpi_bfm_relu3_avmm_0_rw_inst:avs_readdata -> relu3_inst:avmm_0_rw_readdata
	wire  [63:0] relu3_inst_avmm_0_rw_address;                                                                  // relu3_inst:avmm_0_rw_address -> mm_agent_dpi_bfm_relu3_avmm_0_rw_inst:avs_address
	wire   [7:0] relu3_inst_avmm_0_rw_byteenable;                                                               // relu3_inst:avmm_0_rw_byteenable -> mm_agent_dpi_bfm_relu3_avmm_0_rw_inst:avs_byteenable
	wire         relu3_inst_avmm_0_rw_read;                                                                     // relu3_inst:avmm_0_rw_read -> mm_agent_dpi_bfm_relu3_avmm_0_rw_inst:avs_read
	wire         relu3_inst_avmm_0_rw_write;                                                                    // relu3_inst:avmm_0_rw_write -> mm_agent_dpi_bfm_relu3_avmm_0_rw_inst:avs_write
	wire  [63:0] relu3_inst_avmm_0_rw_writedata;                                                                // relu3_inst:avmm_0_rw_writedata -> mm_agent_dpi_bfm_relu3_avmm_0_rw_inst:avs_writedata
	wire  [63:0] relu4_inst_avmm_0_rw_readdata;                                                                 // mm_agent_dpi_bfm_relu4_avmm_0_rw_inst:avs_readdata -> relu4_inst:avmm_0_rw_readdata
	wire  [63:0] relu4_inst_avmm_0_rw_address;                                                                  // relu4_inst:avmm_0_rw_address -> mm_agent_dpi_bfm_relu4_avmm_0_rw_inst:avs_address
	wire   [7:0] relu4_inst_avmm_0_rw_byteenable;                                                               // relu4_inst:avmm_0_rw_byteenable -> mm_agent_dpi_bfm_relu4_avmm_0_rw_inst:avs_byteenable
	wire         relu4_inst_avmm_0_rw_read;                                                                     // relu4_inst:avmm_0_rw_read -> mm_agent_dpi_bfm_relu4_avmm_0_rw_inst:avs_read
	wire         relu4_inst_avmm_0_rw_write;                                                                    // relu4_inst:avmm_0_rw_write -> mm_agent_dpi_bfm_relu4_avmm_0_rw_inst:avs_write
	wire  [63:0] relu4_inst_avmm_0_rw_writedata;                                                                // relu4_inst:avmm_0_rw_writedata -> mm_agent_dpi_bfm_relu4_avmm_0_rw_inst:avs_writedata
	wire  [63:0] softmax_inst_avmm_0_rw_readdata;                                                               // mm_agent_dpi_bfm_softmax_avmm_0_rw_inst:avs_readdata -> softmax_inst:avmm_0_rw_readdata
	wire  [63:0] softmax_inst_avmm_0_rw_address;                                                                // softmax_inst:avmm_0_rw_address -> mm_agent_dpi_bfm_softmax_avmm_0_rw_inst:avs_address
	wire   [7:0] softmax_inst_avmm_0_rw_byteenable;                                                             // softmax_inst:avmm_0_rw_byteenable -> mm_agent_dpi_bfm_softmax_avmm_0_rw_inst:avs_byteenable
	wire         softmax_inst_avmm_0_rw_read;                                                                   // softmax_inst:avmm_0_rw_read -> mm_agent_dpi_bfm_softmax_avmm_0_rw_inst:avs_read
	wire         softmax_inst_avmm_0_rw_write;                                                                  // softmax_inst:avmm_0_rw_write -> mm_agent_dpi_bfm_softmax_avmm_0_rw_inst:avs_write
	wire  [63:0] softmax_inst_avmm_0_rw_writedata;                                                              // softmax_inst:avmm_0_rw_writedata -> mm_agent_dpi_bfm_softmax_avmm_0_rw_inst:avs_writedata
	wire         clock_reset_inst_clock_clk;                                                                    // clock_reset_inst:clock -> [avgpooling1_inst:clock, avgpooling2_inst:clock, component_dpi_controller_avgpooling1_inst:clock, component_dpi_controller_avgpooling2_inst:clock, component_dpi_controller_conv1_inst:clock, component_dpi_controller_conv2_inst:clock, component_dpi_controller_fc1_inst:clock, component_dpi_controller_fc3_inst:clock, component_dpi_controller_relu1_inst:clock, component_dpi_controller_relu2_inst:clock, component_dpi_controller_relu3_inst:clock, component_dpi_controller_relu4_inst:clock, component_dpi_controller_softmax_inst:clock, conv1_inst:clock, conv2_inst:clock, fc1_inst:clock, fc3_inst:clock, irq_mapper:clk, irq_mapper_001:clk, irq_mapper_002:clk, irq_mapper_003:clk, irq_mapper_004:clk, irq_mapper_005:clk, irq_mapper_006:clk, irq_mapper_007:clk, irq_mapper_008:clk, irq_mapper_009:clk, irq_mapper_010:clk, main_dpi_controller_inst:clock, mm_agent_dpi_bfm_avgpooling1_avmm_0_rw_inst:clock, mm_agent_dpi_bfm_avgpooling2_avmm_0_rw_inst:clock, mm_agent_dpi_bfm_conv1_avmm_0_rw_inst:clock, mm_agent_dpi_bfm_conv2_avmm_0_rw_inst:clock, mm_agent_dpi_bfm_fc1_avmm_0_rw_inst:clock, mm_agent_dpi_bfm_fc3_avmm_0_rw_inst:clock, mm_agent_dpi_bfm_relu1_avmm_0_rw_inst:clock, mm_agent_dpi_bfm_relu2_avmm_0_rw_inst:clock, mm_agent_dpi_bfm_relu3_avmm_0_rw_inst:clock, mm_agent_dpi_bfm_relu4_avmm_0_rw_inst:clock, mm_agent_dpi_bfm_softmax_avmm_0_rw_inst:clock, relu1_inst:clock, relu2_inst:clock, relu3_inst:clock, relu4_inst:clock, softmax_inst:clock, stream_source_dpi_bfm_avgpooling1_in0_inst:clock, stream_source_dpi_bfm_avgpooling1_out0_inst:clock, stream_source_dpi_bfm_avgpooling2_in0_inst:clock, stream_source_dpi_bfm_avgpooling2_out0_inst:clock, stream_source_dpi_bfm_conv1_bias_inst:clock, stream_source_dpi_bfm_conv1_in0_inst:clock, stream_source_dpi_bfm_conv1_kernel_inst:clock, stream_source_dpi_bfm_conv1_out0_inst:clock, stream_source_dpi_bfm_conv2_bias_inst:clock, stream_source_dpi_bfm_conv2_in0_inst:clock, stream_source_dpi_bfm_conv2_kernel_inst:clock, stream_source_dpi_bfm_conv2_out0_inst:clock, stream_source_dpi_bfm_fc1_bias_inst:clock, stream_source_dpi_bfm_fc1_in0_inst:clock, stream_source_dpi_bfm_fc1_out0_inst:clock, stream_source_dpi_bfm_fc1_weights_inst:clock, stream_source_dpi_bfm_fc3_bias_inst:clock, stream_source_dpi_bfm_fc3_in0_inst:clock, stream_source_dpi_bfm_fc3_out0_inst:clock, stream_source_dpi_bfm_fc3_weights_inst:clock, stream_source_dpi_bfm_relu1_in0_inst:clock, stream_source_dpi_bfm_relu1_out0_inst:clock, stream_source_dpi_bfm_relu2_in0_inst:clock, stream_source_dpi_bfm_relu2_out0_inst:clock, stream_source_dpi_bfm_relu3_in0_inst:clock, stream_source_dpi_bfm_relu3_out0_inst:clock, stream_source_dpi_bfm_relu4_in0_inst:clock, stream_source_dpi_bfm_relu4_out0_inst:clock, stream_source_dpi_bfm_softmax_in0_inst:clock, stream_source_dpi_bfm_softmax_out0_inst:clock]
	wire         clock_reset_inst_clock2x_clk;                                                                  // clock_reset_inst:clock2x -> [component_dpi_controller_avgpooling1_inst:clock2x, component_dpi_controller_avgpooling2_inst:clock2x, component_dpi_controller_conv1_inst:clock2x, component_dpi_controller_conv2_inst:clock2x, component_dpi_controller_fc1_inst:clock2x, component_dpi_controller_fc3_inst:clock2x, component_dpi_controller_relu1_inst:clock2x, component_dpi_controller_relu2_inst:clock2x, component_dpi_controller_relu3_inst:clock2x, component_dpi_controller_relu4_inst:clock2x, component_dpi_controller_softmax_inst:clock2x, main_dpi_controller_inst:clock2x, stream_source_dpi_bfm_avgpooling1_in0_inst:clock2x, stream_source_dpi_bfm_avgpooling1_out0_inst:clock2x, stream_source_dpi_bfm_avgpooling2_in0_inst:clock2x, stream_source_dpi_bfm_avgpooling2_out0_inst:clock2x, stream_source_dpi_bfm_conv1_bias_inst:clock2x, stream_source_dpi_bfm_conv1_in0_inst:clock2x, stream_source_dpi_bfm_conv1_kernel_inst:clock2x, stream_source_dpi_bfm_conv1_out0_inst:clock2x, stream_source_dpi_bfm_conv2_bias_inst:clock2x, stream_source_dpi_bfm_conv2_in0_inst:clock2x, stream_source_dpi_bfm_conv2_kernel_inst:clock2x, stream_source_dpi_bfm_conv2_out0_inst:clock2x, stream_source_dpi_bfm_fc1_bias_inst:clock2x, stream_source_dpi_bfm_fc1_in0_inst:clock2x, stream_source_dpi_bfm_fc1_out0_inst:clock2x, stream_source_dpi_bfm_fc1_weights_inst:clock2x, stream_source_dpi_bfm_fc3_bias_inst:clock2x, stream_source_dpi_bfm_fc3_in0_inst:clock2x, stream_source_dpi_bfm_fc3_out0_inst:clock2x, stream_source_dpi_bfm_fc3_weights_inst:clock2x, stream_source_dpi_bfm_relu1_in0_inst:clock2x, stream_source_dpi_bfm_relu1_out0_inst:clock2x, stream_source_dpi_bfm_relu2_in0_inst:clock2x, stream_source_dpi_bfm_relu2_out0_inst:clock2x, stream_source_dpi_bfm_relu3_in0_inst:clock2x, stream_source_dpi_bfm_relu3_out0_inst:clock2x, stream_source_dpi_bfm_relu4_in0_inst:clock2x, stream_source_dpi_bfm_relu4_out0_inst:clock2x, stream_source_dpi_bfm_softmax_in0_inst:clock2x, stream_source_dpi_bfm_softmax_out0_inst:clock2x]
	wire         component_dpi_controller_avgpooling1_inst_component_call_valid;                                // component_dpi_controller_avgpooling1_inst:start -> avgpooling1_inst:start
	wire         avgpooling1_inst_call_stall;                                                                   // avgpooling1_inst:busy -> component_dpi_controller_avgpooling1_inst:busy
	wire         component_dpi_controller_avgpooling2_inst_component_call_valid;                                // component_dpi_controller_avgpooling2_inst:start -> avgpooling2_inst:start
	wire         avgpooling2_inst_call_stall;                                                                   // avgpooling2_inst:busy -> component_dpi_controller_avgpooling2_inst:busy
	wire         component_dpi_controller_conv1_inst_component_call_valid;                                      // component_dpi_controller_conv1_inst:start -> conv1_inst:start
	wire         conv1_inst_call_stall;                                                                         // conv1_inst:busy -> component_dpi_controller_conv1_inst:busy
	wire         component_dpi_controller_conv2_inst_component_call_valid;                                      // component_dpi_controller_conv2_inst:start -> conv2_inst:start
	wire         conv2_inst_call_stall;                                                                         // conv2_inst:busy -> component_dpi_controller_conv2_inst:busy
	wire         component_dpi_controller_fc1_inst_component_call_valid;                                        // component_dpi_controller_fc1_inst:start -> fc1_inst:start
	wire         fc1_inst_call_stall;                                                                           // fc1_inst:busy -> component_dpi_controller_fc1_inst:busy
	wire         component_dpi_controller_fc3_inst_component_call_valid;                                        // component_dpi_controller_fc3_inst:start -> fc3_inst:start
	wire         fc3_inst_call_stall;                                                                           // fc3_inst:busy -> component_dpi_controller_fc3_inst:busy
	wire         component_dpi_controller_relu1_inst_component_call_valid;                                      // component_dpi_controller_relu1_inst:start -> relu1_inst:start
	wire         relu1_inst_call_stall;                                                                         // relu1_inst:busy -> component_dpi_controller_relu1_inst:busy
	wire         component_dpi_controller_relu2_inst_component_call_valid;                                      // component_dpi_controller_relu2_inst:start -> relu2_inst:start
	wire         relu2_inst_call_stall;                                                                         // relu2_inst:busy -> component_dpi_controller_relu2_inst:busy
	wire         component_dpi_controller_relu3_inst_component_call_valid;                                      // component_dpi_controller_relu3_inst:start -> relu3_inst:start
	wire         relu3_inst_call_stall;                                                                         // relu3_inst:busy -> component_dpi_controller_relu3_inst:busy
	wire         component_dpi_controller_relu4_inst_component_call_valid;                                      // component_dpi_controller_relu4_inst:start -> relu4_inst:start
	wire         relu4_inst_call_stall;                                                                         // relu4_inst:busy -> component_dpi_controller_relu4_inst:busy
	wire         component_dpi_controller_softmax_inst_component_call_valid;                                    // component_dpi_controller_softmax_inst:start -> softmax_inst:start
	wire         softmax_inst_call_stall;                                                                       // softmax_inst:busy -> component_dpi_controller_softmax_inst:busy
	wire         component_dpi_controller_avgpooling1_inst_component_done_conduit;                              // component_dpi_controller_avgpooling1_inst:component_done -> concatenate_component_done_inst:in_conduit_0
	wire         component_dpi_controller_avgpooling2_inst_component_done_conduit;                              // component_dpi_controller_avgpooling2_inst:component_done -> concatenate_component_done_inst:in_conduit_1
	wire         component_dpi_controller_softmax_inst_component_done_conduit;                                  // component_dpi_controller_softmax_inst:component_done -> concatenate_component_done_inst:in_conduit_10
	wire         component_dpi_controller_conv1_inst_component_done_conduit;                                    // component_dpi_controller_conv1_inst:component_done -> concatenate_component_done_inst:in_conduit_2
	wire         component_dpi_controller_conv2_inst_component_done_conduit;                                    // component_dpi_controller_conv2_inst:component_done -> concatenate_component_done_inst:in_conduit_3
	wire         component_dpi_controller_fc1_inst_component_done_conduit;                                      // component_dpi_controller_fc1_inst:component_done -> concatenate_component_done_inst:in_conduit_4
	wire         component_dpi_controller_fc3_inst_component_done_conduit;                                      // component_dpi_controller_fc3_inst:component_done -> concatenate_component_done_inst:in_conduit_5
	wire         component_dpi_controller_relu1_inst_component_done_conduit;                                    // component_dpi_controller_relu1_inst:component_done -> concatenate_component_done_inst:in_conduit_6
	wire         component_dpi_controller_relu2_inst_component_done_conduit;                                    // component_dpi_controller_relu2_inst:component_done -> concatenate_component_done_inst:in_conduit_7
	wire         component_dpi_controller_relu3_inst_component_done_conduit;                                    // component_dpi_controller_relu3_inst:component_done -> concatenate_component_done_inst:in_conduit_8
	wire         component_dpi_controller_relu4_inst_component_done_conduit;                                    // component_dpi_controller_relu4_inst:component_done -> concatenate_component_done_inst:in_conduit_9
	wire  [10:0] main_dpi_controller_inst_component_enabled_conduit;                                            // main_dpi_controller_inst:component_enabled -> split_component_start_inst:in_conduit
	wire         component_dpi_controller_avgpooling1_inst_component_wait_for_stream_writes_conduit;            // component_dpi_controller_avgpooling1_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_0
	wire         component_dpi_controller_avgpooling2_inst_component_wait_for_stream_writes_conduit;            // component_dpi_controller_avgpooling2_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_1
	wire         component_dpi_controller_softmax_inst_component_wait_for_stream_writes_conduit;                // component_dpi_controller_softmax_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_10
	wire         component_dpi_controller_conv1_inst_component_wait_for_stream_writes_conduit;                  // component_dpi_controller_conv1_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_2
	wire         component_dpi_controller_conv2_inst_component_wait_for_stream_writes_conduit;                  // component_dpi_controller_conv2_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_3
	wire         component_dpi_controller_fc1_inst_component_wait_for_stream_writes_conduit;                    // component_dpi_controller_fc1_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_4
	wire         component_dpi_controller_fc3_inst_component_wait_for_stream_writes_conduit;                    // component_dpi_controller_fc3_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_5
	wire         component_dpi_controller_relu1_inst_component_wait_for_stream_writes_conduit;                  // component_dpi_controller_relu1_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_6
	wire         component_dpi_controller_relu2_inst_component_wait_for_stream_writes_conduit;                  // component_dpi_controller_relu2_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_7
	wire         component_dpi_controller_relu3_inst_component_wait_for_stream_writes_conduit;                  // component_dpi_controller_relu3_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_8
	wire         component_dpi_controller_relu4_inst_component_wait_for_stream_writes_conduit;                  // component_dpi_controller_relu4_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_9
	wire         component_dpi_controller_avgpooling1_inst_dpi_control_bind_conduit;                            // component_dpi_controller_avgpooling1_inst:bind_interfaces -> avgpooling1_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_avgpooling2_inst_dpi_control_bind_conduit;                            // component_dpi_controller_avgpooling2_inst:bind_interfaces -> avgpooling2_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_conv1_inst_dpi_control_bind_conduit;                                  // component_dpi_controller_conv1_inst:bind_interfaces -> conv1_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_conv2_inst_dpi_control_bind_conduit;                                  // component_dpi_controller_conv2_inst:bind_interfaces -> conv2_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_fc1_inst_dpi_control_bind_conduit;                                    // component_dpi_controller_fc1_inst:bind_interfaces -> fc1_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_fc3_inst_dpi_control_bind_conduit;                                    // component_dpi_controller_fc3_inst:bind_interfaces -> fc3_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_relu1_inst_dpi_control_bind_conduit;                                  // component_dpi_controller_relu1_inst:bind_interfaces -> relu1_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_relu2_inst_dpi_control_bind_conduit;                                  // component_dpi_controller_relu2_inst:bind_interfaces -> relu2_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_relu3_inst_dpi_control_bind_conduit;                                  // component_dpi_controller_relu3_inst:bind_interfaces -> relu3_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_relu4_inst_dpi_control_bind_conduit;                                  // component_dpi_controller_relu4_inst:bind_interfaces -> relu4_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_softmax_inst_dpi_control_bind_conduit;                                // component_dpi_controller_softmax_inst:bind_interfaces -> softmax_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_avgpooling1_inst_dpi_control_enable_conduit;                          // component_dpi_controller_avgpooling1_inst:enable_interfaces -> avgpooling1_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_avgpooling2_inst_dpi_control_enable_conduit;                          // component_dpi_controller_avgpooling2_inst:enable_interfaces -> avgpooling2_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_conv1_inst_dpi_control_enable_conduit;                                // component_dpi_controller_conv1_inst:enable_interfaces -> conv1_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_conv2_inst_dpi_control_enable_conduit;                                // component_dpi_controller_conv2_inst:enable_interfaces -> conv2_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_fc1_inst_dpi_control_enable_conduit;                                  // component_dpi_controller_fc1_inst:enable_interfaces -> fc1_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_fc3_inst_dpi_control_enable_conduit;                                  // component_dpi_controller_fc3_inst:enable_interfaces -> fc3_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_relu1_inst_dpi_control_enable_conduit;                                // component_dpi_controller_relu1_inst:enable_interfaces -> relu1_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_relu2_inst_dpi_control_enable_conduit;                                // component_dpi_controller_relu2_inst:enable_interfaces -> relu2_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_relu3_inst_dpi_control_enable_conduit;                                // component_dpi_controller_relu3_inst:enable_interfaces -> relu3_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_relu4_inst_dpi_control_enable_conduit;                                // component_dpi_controller_relu4_inst:enable_interfaces -> relu4_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_softmax_inst_dpi_control_enable_conduit;                              // component_dpi_controller_softmax_inst:enable_interfaces -> softmax_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire  [10:0] concatenate_component_done_inst_out_conduit_conduit;                                           // concatenate_component_done_inst:out_conduit -> main_dpi_controller_inst:component_done
	wire  [10:0] concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit;                         // concatenate_component_wait_for_stream_writes_inst:out_conduit -> main_dpi_controller_inst:component_wait_for_stream_writes
	wire         split_component_start_inst_out_conduit_0_conduit;                                              // split_component_start_inst:out_conduit_0 -> component_dpi_controller_avgpooling1_inst:component_enabled
	wire         avgpooling1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;           // avgpooling1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_avgpooling1_avmm_0_rw_inst:do_bind
	wire         avgpooling2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;           // avgpooling2_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_avgpooling2_avmm_0_rw_inst:do_bind
	wire         conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;                 // conv1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_conv1_avmm_0_rw_inst:do_bind
	wire         conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;                 // conv2_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_conv2_avmm_0_rw_inst:do_bind
	wire         fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;                   // fc1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_fc1_avmm_0_rw_inst:do_bind
	wire         fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;                   // fc3_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_fc3_avmm_0_rw_inst:do_bind
	wire         relu1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;                 // relu1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_relu1_avmm_0_rw_inst:do_bind
	wire         relu2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;                 // relu2_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_relu2_avmm_0_rw_inst:do_bind
	wire         relu3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;                 // relu3_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_relu3_avmm_0_rw_inst:do_bind
	wire         relu4_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;                 // relu4_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_relu4_avmm_0_rw_inst:do_bind
	wire         softmax_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;               // softmax_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_softmax_avmm_0_rw_inst:do_bind
	wire         avgpooling1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;         // avgpooling1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_avgpooling1_avmm_0_rw_inst:enable
	wire         avgpooling2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;         // avgpooling2_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_avgpooling2_avmm_0_rw_inst:enable
	wire         conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;               // conv1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_conv1_avmm_0_rw_inst:enable
	wire         conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;               // conv2_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_conv2_avmm_0_rw_inst:enable
	wire         fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;                 // fc1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_fc1_avmm_0_rw_inst:enable
	wire         fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;                 // fc3_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_fc3_avmm_0_rw_inst:enable
	wire         relu1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;               // relu1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_relu1_avmm_0_rw_inst:enable
	wire         relu2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;               // relu2_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_relu2_avmm_0_rw_inst:enable
	wire         relu3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;               // relu3_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_relu3_avmm_0_rw_inst:enable
	wire         relu4_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;               // relu4_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_relu4_avmm_0_rw_inst:enable
	wire         softmax_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;             // softmax_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> mm_agent_dpi_bfm_softmax_avmm_0_rw_inst:enable
	wire         avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit; // avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_avgpooling1_in0_inst:source_ready
	wire         avgpooling2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit; // avgpooling2_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_avgpooling2_in0_inst:source_ready
	wire         conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit;       // conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_conv1_bias_inst:source_ready
	wire         conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit;       // conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_conv2_bias_inst:source_ready
	wire         fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit;         // fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_fc1_bias_inst:source_ready
	wire         fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit;         // fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_fc3_bias_inst:source_ready
	wire         relu1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit;       // relu1_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_relu1_in0_inst:source_ready
	wire         relu2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit;       // relu2_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_relu2_in0_inst:source_ready
	wire         relu3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit;       // relu3_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_relu3_in0_inst:source_ready
	wire         relu4_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit;       // relu4_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_relu4_in0_inst:source_ready
	wire         softmax_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit;     // softmax_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_softmax_in0_inst:source_ready
	wire         split_component_start_inst_out_conduit_1_conduit;                                              // split_component_start_inst:out_conduit_1 -> component_dpi_controller_avgpooling2_inst:component_enabled
	wire         avgpooling1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;           // avgpooling1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_avgpooling1_in0_inst:do_bind
	wire         avgpooling2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;           // avgpooling2_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_avgpooling2_in0_inst:do_bind
	wire         conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;                 // conv1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_conv1_bias_inst:do_bind
	wire         conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;                 // conv2_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_conv2_bias_inst:do_bind
	wire         fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;                   // fc1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_fc1_bias_inst:do_bind
	wire         fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;                   // fc3_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_fc3_bias_inst:do_bind
	wire         relu1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;                 // relu1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_relu1_in0_inst:do_bind
	wire         relu2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;                 // relu2_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_relu2_in0_inst:do_bind
	wire         relu3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;                 // relu3_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_relu3_in0_inst:do_bind
	wire         relu4_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;                 // relu4_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_relu4_in0_inst:do_bind
	wire         softmax_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;               // softmax_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_softmax_in0_inst:do_bind
	wire         avgpooling1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;         // avgpooling1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_avgpooling1_in0_inst:enable
	wire         avgpooling2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;         // avgpooling2_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_avgpooling2_in0_inst:enable
	wire         conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;               // conv1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_conv1_bias_inst:enable
	wire         conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;               // conv2_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_conv2_bias_inst:enable
	wire         fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;                 // fc1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_fc1_bias_inst:enable
	wire         fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;                 // fc3_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_fc3_bias_inst:enable
	wire         relu1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;               // relu1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_relu1_in0_inst:enable
	wire         relu2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;               // relu2_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_relu2_in0_inst:enable
	wire         relu3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;               // relu3_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_relu3_in0_inst:enable
	wire         relu4_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;               // relu4_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_relu4_in0_inst:enable
	wire         softmax_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;             // softmax_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_softmax_in0_inst:enable
	wire         avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit; // avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_avgpooling1_out0_inst:source_ready
	wire         avgpooling2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit; // avgpooling2_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_avgpooling2_out0_inst:source_ready
	wire         conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit;       // conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_conv1_in0_inst:source_ready
	wire         conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit;       // conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_conv2_in0_inst:source_ready
	wire         fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit;         // fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_fc1_in0_inst:source_ready
	wire         fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit;         // fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_fc3_in0_inst:source_ready
	wire         relu1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit;       // relu1_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_relu1_out0_inst:source_ready
	wire         relu2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit;       // relu2_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_relu2_out0_inst:source_ready
	wire         relu3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit;       // relu3_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_relu3_out0_inst:source_ready
	wire         relu4_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit;       // relu4_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_relu4_out0_inst:source_ready
	wire         softmax_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit;     // softmax_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_softmax_out0_inst:source_ready
	wire         split_component_start_inst_out_conduit_10_conduit;                                             // split_component_start_inst:out_conduit_10 -> component_dpi_controller_softmax_inst:component_enabled
	wire         split_component_start_inst_out_conduit_2_conduit;                                              // split_component_start_inst:out_conduit_2 -> component_dpi_controller_conv1_inst:component_enabled
	wire         avgpooling1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;           // avgpooling1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_avgpooling1_out0_inst:do_bind
	wire         avgpooling2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;           // avgpooling2_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_avgpooling2_out0_inst:do_bind
	wire         conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;                 // conv1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_conv1_in0_inst:do_bind
	wire         conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;                 // conv2_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_conv2_in0_inst:do_bind
	wire         fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;                   // fc1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_fc1_in0_inst:do_bind
	wire         fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;                   // fc3_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_fc3_in0_inst:do_bind
	wire         relu1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;                 // relu1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_relu1_out0_inst:do_bind
	wire         relu2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;                 // relu2_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_relu2_out0_inst:do_bind
	wire         relu3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;                 // relu3_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_relu3_out0_inst:do_bind
	wire         relu4_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;                 // relu4_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_relu4_out0_inst:do_bind
	wire         softmax_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;               // softmax_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_softmax_out0_inst:do_bind
	wire         avgpooling1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;         // avgpooling1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_avgpooling1_out0_inst:enable
	wire         avgpooling2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;         // avgpooling2_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_avgpooling2_out0_inst:enable
	wire         conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;               // conv1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_conv1_in0_inst:enable
	wire         conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;               // conv2_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_conv2_in0_inst:enable
	wire         fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;                 // fc1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_fc1_in0_inst:enable
	wire         fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;                 // fc3_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_fc3_in0_inst:enable
	wire         relu1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;               // relu1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_relu1_out0_inst:enable
	wire         relu2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;               // relu2_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_relu2_out0_inst:enable
	wire         relu3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;               // relu3_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_relu3_out0_inst:enable
	wire         relu4_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;               // relu4_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_relu4_out0_inst:enable
	wire         softmax_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;             // softmax_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_softmax_out0_inst:enable
	wire         conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit;       // conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_conv1_kernel_inst:source_ready
	wire         conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit;       // conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_conv2_kernel_inst:source_ready
	wire         fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit;         // fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_fc1_out0_inst:source_ready
	wire         fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit;         // fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_fc3_out0_inst:source_ready
	wire         split_component_start_inst_out_conduit_3_conduit;                                              // split_component_start_inst:out_conduit_3 -> component_dpi_controller_conv2_inst:component_enabled
	wire         conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit;                 // conv1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_conv1_kernel_inst:do_bind
	wire         conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit;                 // conv2_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_conv2_kernel_inst:do_bind
	wire         fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit;                   // fc1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_fc1_out0_inst:do_bind
	wire         fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit;                   // fc3_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_fc3_out0_inst:do_bind
	wire         conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit;               // conv1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_conv1_kernel_inst:enable
	wire         conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit;               // conv2_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_conv2_kernel_inst:enable
	wire         fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit;                 // fc1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_fc1_out0_inst:enable
	wire         fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit;                 // fc3_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_fc3_out0_inst:enable
	wire         conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit;       // conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_conv1_out0_inst:source_ready
	wire         conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit;       // conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_conv2_out0_inst:source_ready
	wire         fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit;         // fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_fc1_weights_inst:source_ready
	wire         fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit;         // fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_fc3_weights_inst:source_ready
	wire         split_component_start_inst_out_conduit_4_conduit;                                              // split_component_start_inst:out_conduit_4 -> component_dpi_controller_fc1_inst:component_enabled
	wire         conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit;                 // conv1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_conv1_out0_inst:do_bind
	wire         conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit;                 // conv2_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_conv2_out0_inst:do_bind
	wire         fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit;                   // fc1_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_fc1_weights_inst:do_bind
	wire         fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit;                   // fc3_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_fc3_weights_inst:do_bind
	wire         conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit;               // conv1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_conv1_out0_inst:enable
	wire         conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit;               // conv2_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_conv2_out0_inst:enable
	wire         fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit;                 // fc1_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_fc1_weights_inst:enable
	wire         fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit;                 // fc3_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_fc3_weights_inst:enable
	wire         split_component_start_inst_out_conduit_5_conduit;                                              // split_component_start_inst:out_conduit_5 -> component_dpi_controller_fc3_inst:component_enabled
	wire         split_component_start_inst_out_conduit_6_conduit;                                              // split_component_start_inst:out_conduit_6 -> component_dpi_controller_relu1_inst:component_enabled
	wire         split_component_start_inst_out_conduit_7_conduit;                                              // split_component_start_inst:out_conduit_7 -> component_dpi_controller_relu2_inst:component_enabled
	wire         split_component_start_inst_out_conduit_8_conduit;                                              // split_component_start_inst:out_conduit_8 -> component_dpi_controller_relu3_inst:component_enabled
	wire         split_component_start_inst_out_conduit_9_conduit;                                              // split_component_start_inst:out_conduit_9 -> component_dpi_controller_relu4_inst:component_enabled
	wire         component_dpi_controller_avgpooling1_inst_read_implicit_streams_conduit;                       // component_dpi_controller_avgpooling1_inst:read_implicit_streams -> avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_avgpooling2_inst_read_implicit_streams_conduit;                       // component_dpi_controller_avgpooling2_inst:read_implicit_streams -> avgpooling2_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_conv1_inst_read_implicit_streams_conduit;                             // component_dpi_controller_conv1_inst:read_implicit_streams -> conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_conv2_inst_read_implicit_streams_conduit;                             // component_dpi_controller_conv2_inst:read_implicit_streams -> conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_fc1_inst_read_implicit_streams_conduit;                               // component_dpi_controller_fc1_inst:read_implicit_streams -> fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_fc3_inst_read_implicit_streams_conduit;                               // component_dpi_controller_fc3_inst:read_implicit_streams -> fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_relu1_inst_read_implicit_streams_conduit;                             // component_dpi_controller_relu1_inst:read_implicit_streams -> relu1_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_relu2_inst_read_implicit_streams_conduit;                             // component_dpi_controller_relu2_inst:read_implicit_streams -> relu2_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_relu3_inst_read_implicit_streams_conduit;                             // component_dpi_controller_relu3_inst:read_implicit_streams -> relu3_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_relu4_inst_read_implicit_streams_conduit;                             // component_dpi_controller_relu4_inst:read_implicit_streams -> relu4_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_softmax_inst_read_implicit_streams_conduit;                           // component_dpi_controller_softmax_inst:read_implicit_streams -> softmax_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         main_dpi_controller_inst_reset_ctrl_conduit;                                                   // main_dpi_controller_inst:trigger_reset -> clock_reset_inst:trigger_reset
	wire         avgpooling1_inst_return_valid;                                                                 // avgpooling1_inst:done -> component_dpi_controller_avgpooling1_inst:done
	wire         component_dpi_controller_avgpooling1_inst_component_return_stall;                              // component_dpi_controller_avgpooling1_inst:stall -> avgpooling1_inst:stall
	wire         avgpooling2_inst_return_valid;                                                                 // avgpooling2_inst:done -> component_dpi_controller_avgpooling2_inst:done
	wire         component_dpi_controller_avgpooling2_inst_component_return_stall;                              // component_dpi_controller_avgpooling2_inst:stall -> avgpooling2_inst:stall
	wire         conv1_inst_return_valid;                                                                       // conv1_inst:done -> component_dpi_controller_conv1_inst:done
	wire         component_dpi_controller_conv1_inst_component_return_stall;                                    // component_dpi_controller_conv1_inst:stall -> conv1_inst:stall
	wire         conv2_inst_return_valid;                                                                       // conv2_inst:done -> component_dpi_controller_conv2_inst:done
	wire         component_dpi_controller_conv2_inst_component_return_stall;                                    // component_dpi_controller_conv2_inst:stall -> conv2_inst:stall
	wire         fc1_inst_return_valid;                                                                         // fc1_inst:done -> component_dpi_controller_fc1_inst:done
	wire         component_dpi_controller_fc1_inst_component_return_stall;                                      // component_dpi_controller_fc1_inst:stall -> fc1_inst:stall
	wire         fc3_inst_return_valid;                                                                         // fc3_inst:done -> component_dpi_controller_fc3_inst:done
	wire         component_dpi_controller_fc3_inst_component_return_stall;                                      // component_dpi_controller_fc3_inst:stall -> fc3_inst:stall
	wire         relu1_inst_return_valid;                                                                       // relu1_inst:done -> component_dpi_controller_relu1_inst:done
	wire         component_dpi_controller_relu1_inst_component_return_stall;                                    // component_dpi_controller_relu1_inst:stall -> relu1_inst:stall
	wire         relu2_inst_return_valid;                                                                       // relu2_inst:done -> component_dpi_controller_relu2_inst:done
	wire         component_dpi_controller_relu2_inst_component_return_stall;                                    // component_dpi_controller_relu2_inst:stall -> relu2_inst:stall
	wire         relu3_inst_return_valid;                                                                       // relu3_inst:done -> component_dpi_controller_relu3_inst:done
	wire         component_dpi_controller_relu3_inst_component_return_stall;                                    // component_dpi_controller_relu3_inst:stall -> relu3_inst:stall
	wire         relu4_inst_return_valid;                                                                       // relu4_inst:done -> component_dpi_controller_relu4_inst:done
	wire         component_dpi_controller_relu4_inst_component_return_stall;                                    // component_dpi_controller_relu4_inst:stall -> relu4_inst:stall
	wire         softmax_inst_return_valid;                                                                     // softmax_inst:done -> component_dpi_controller_softmax_inst:done
	wire         component_dpi_controller_softmax_inst_component_return_stall;                                  // component_dpi_controller_softmax_inst:stall -> softmax_inst:stall
	wire  [63:0] stream_source_dpi_bfm_conv1_bias_inst_source_data_data;                                        // stream_source_dpi_bfm_conv1_bias_inst:source_data -> conv1_inst:bias
	wire  [63:0] stream_source_dpi_bfm_conv2_bias_inst_source_data_data;                                        // stream_source_dpi_bfm_conv2_bias_inst:source_data -> conv2_inst:bias
	wire  [63:0] stream_source_dpi_bfm_fc1_bias_inst_source_data_data;                                          // stream_source_dpi_bfm_fc1_bias_inst:source_data -> fc1_inst:bias
	wire  [63:0] stream_source_dpi_bfm_fc3_bias_inst_source_data_data;                                          // stream_source_dpi_bfm_fc3_bias_inst:source_data -> fc3_inst:bias
	wire  [63:0] stream_source_dpi_bfm_avgpooling1_in0_inst_source_data_data;                                   // stream_source_dpi_bfm_avgpooling1_in0_inst:source_data -> avgpooling1_inst:in0
	wire  [63:0] stream_source_dpi_bfm_avgpooling2_in0_inst_source_data_data;                                   // stream_source_dpi_bfm_avgpooling2_in0_inst:source_data -> avgpooling2_inst:in0
	wire  [63:0] stream_source_dpi_bfm_conv1_in0_inst_source_data_data;                                         // stream_source_dpi_bfm_conv1_in0_inst:source_data -> conv1_inst:in0
	wire  [63:0] stream_source_dpi_bfm_conv2_in0_inst_source_data_data;                                         // stream_source_dpi_bfm_conv2_in0_inst:source_data -> conv2_inst:in0
	wire  [63:0] stream_source_dpi_bfm_fc1_in0_inst_source_data_data;                                           // stream_source_dpi_bfm_fc1_in0_inst:source_data -> fc1_inst:in0
	wire  [63:0] stream_source_dpi_bfm_fc3_in0_inst_source_data_data;                                           // stream_source_dpi_bfm_fc3_in0_inst:source_data -> fc3_inst:in0
	wire  [63:0] stream_source_dpi_bfm_relu1_in0_inst_source_data_data;                                         // stream_source_dpi_bfm_relu1_in0_inst:source_data -> relu1_inst:in0
	wire  [63:0] stream_source_dpi_bfm_relu2_in0_inst_source_data_data;                                         // stream_source_dpi_bfm_relu2_in0_inst:source_data -> relu2_inst:in0
	wire  [63:0] stream_source_dpi_bfm_relu3_in0_inst_source_data_data;                                         // stream_source_dpi_bfm_relu3_in0_inst:source_data -> relu3_inst:in0
	wire  [63:0] stream_source_dpi_bfm_relu4_in0_inst_source_data_data;                                         // stream_source_dpi_bfm_relu4_in0_inst:source_data -> relu4_inst:in0
	wire  [63:0] stream_source_dpi_bfm_softmax_in0_inst_source_data_data;                                       // stream_source_dpi_bfm_softmax_in0_inst:source_data -> softmax_inst:in0
	wire  [63:0] stream_source_dpi_bfm_conv1_kernel_inst_source_data_data;                                      // stream_source_dpi_bfm_conv1_kernel_inst:source_data -> conv1_inst:kernel
	wire  [63:0] stream_source_dpi_bfm_conv2_kernel_inst_source_data_data;                                      // stream_source_dpi_bfm_conv2_kernel_inst:source_data -> conv2_inst:kernel
	wire  [63:0] stream_source_dpi_bfm_avgpooling1_out0_inst_source_data_data;                                  // stream_source_dpi_bfm_avgpooling1_out0_inst:source_data -> avgpooling1_inst:out0
	wire  [63:0] stream_source_dpi_bfm_avgpooling2_out0_inst_source_data_data;                                  // stream_source_dpi_bfm_avgpooling2_out0_inst:source_data -> avgpooling2_inst:out0
	wire  [63:0] stream_source_dpi_bfm_conv1_out0_inst_source_data_data;                                        // stream_source_dpi_bfm_conv1_out0_inst:source_data -> conv1_inst:out0
	wire  [63:0] stream_source_dpi_bfm_conv2_out0_inst_source_data_data;                                        // stream_source_dpi_bfm_conv2_out0_inst:source_data -> conv2_inst:out0
	wire  [63:0] stream_source_dpi_bfm_fc1_out0_inst_source_data_data;                                          // stream_source_dpi_bfm_fc1_out0_inst:source_data -> fc1_inst:out0
	wire  [63:0] stream_source_dpi_bfm_fc3_out0_inst_source_data_data;                                          // stream_source_dpi_bfm_fc3_out0_inst:source_data -> fc3_inst:out0
	wire  [63:0] stream_source_dpi_bfm_relu1_out0_inst_source_data_data;                                        // stream_source_dpi_bfm_relu1_out0_inst:source_data -> relu1_inst:out0
	wire  [63:0] stream_source_dpi_bfm_relu2_out0_inst_source_data_data;                                        // stream_source_dpi_bfm_relu2_out0_inst:source_data -> relu2_inst:out0
	wire  [63:0] stream_source_dpi_bfm_relu3_out0_inst_source_data_data;                                        // stream_source_dpi_bfm_relu3_out0_inst:source_data -> relu3_inst:out0
	wire  [63:0] stream_source_dpi_bfm_relu4_out0_inst_source_data_data;                                        // stream_source_dpi_bfm_relu4_out0_inst:source_data -> relu4_inst:out0
	wire  [63:0] stream_source_dpi_bfm_softmax_out0_inst_source_data_data;                                      // stream_source_dpi_bfm_softmax_out0_inst:source_data -> softmax_inst:out0
	wire  [63:0] stream_source_dpi_bfm_fc1_weights_inst_source_data_data;                                       // stream_source_dpi_bfm_fc1_weights_inst:source_data -> fc1_inst:weights
	wire  [63:0] stream_source_dpi_bfm_fc3_weights_inst_source_data_data;                                       // stream_source_dpi_bfm_fc3_weights_inst:source_data -> fc3_inst:weights
	wire         clock_reset_inst_reset_reset;                                                                  // clock_reset_inst:resetn -> [avgpooling1_inst:resetn, avgpooling2_inst:resetn, component_dpi_controller_avgpooling1_inst:resetn, component_dpi_controller_avgpooling2_inst:resetn, component_dpi_controller_conv1_inst:resetn, component_dpi_controller_conv2_inst:resetn, component_dpi_controller_fc1_inst:resetn, component_dpi_controller_fc3_inst:resetn, component_dpi_controller_relu1_inst:resetn, component_dpi_controller_relu2_inst:resetn, component_dpi_controller_relu3_inst:resetn, component_dpi_controller_relu4_inst:resetn, component_dpi_controller_softmax_inst:resetn, conv1_inst:resetn, conv2_inst:resetn, fc1_inst:resetn, fc3_inst:resetn, irq_mapper:reset, irq_mapper_001:reset, irq_mapper_002:reset, irq_mapper_003:reset, irq_mapper_004:reset, irq_mapper_005:reset, irq_mapper_006:reset, irq_mapper_007:reset, irq_mapper_008:reset, irq_mapper_009:reset, irq_mapper_010:reset, main_dpi_controller_inst:resetn, mm_agent_dpi_bfm_avgpooling1_avmm_0_rw_inst:reset_n, mm_agent_dpi_bfm_avgpooling2_avmm_0_rw_inst:reset_n, mm_agent_dpi_bfm_conv1_avmm_0_rw_inst:reset_n, mm_agent_dpi_bfm_conv2_avmm_0_rw_inst:reset_n, mm_agent_dpi_bfm_fc1_avmm_0_rw_inst:reset_n, mm_agent_dpi_bfm_fc3_avmm_0_rw_inst:reset_n, mm_agent_dpi_bfm_relu1_avmm_0_rw_inst:reset_n, mm_agent_dpi_bfm_relu2_avmm_0_rw_inst:reset_n, mm_agent_dpi_bfm_relu3_avmm_0_rw_inst:reset_n, mm_agent_dpi_bfm_relu4_avmm_0_rw_inst:reset_n, mm_agent_dpi_bfm_softmax_avmm_0_rw_inst:reset_n, relu1_inst:resetn, relu2_inst:resetn, relu3_inst:resetn, relu4_inst:resetn, softmax_inst:resetn, stream_source_dpi_bfm_avgpooling1_in0_inst:resetn, stream_source_dpi_bfm_avgpooling1_out0_inst:resetn, stream_source_dpi_bfm_avgpooling2_in0_inst:resetn, stream_source_dpi_bfm_avgpooling2_out0_inst:resetn, stream_source_dpi_bfm_conv1_bias_inst:resetn, stream_source_dpi_bfm_conv1_in0_inst:resetn, stream_source_dpi_bfm_conv1_kernel_inst:resetn, stream_source_dpi_bfm_conv1_out0_inst:resetn, stream_source_dpi_bfm_conv2_bias_inst:resetn, stream_source_dpi_bfm_conv2_in0_inst:resetn, stream_source_dpi_bfm_conv2_kernel_inst:resetn, stream_source_dpi_bfm_conv2_out0_inst:resetn, stream_source_dpi_bfm_fc1_bias_inst:resetn, stream_source_dpi_bfm_fc1_in0_inst:resetn, stream_source_dpi_bfm_fc1_out0_inst:resetn, stream_source_dpi_bfm_fc1_weights_inst:resetn, stream_source_dpi_bfm_fc3_bias_inst:resetn, stream_source_dpi_bfm_fc3_in0_inst:resetn, stream_source_dpi_bfm_fc3_out0_inst:resetn, stream_source_dpi_bfm_fc3_weights_inst:resetn, stream_source_dpi_bfm_relu1_in0_inst:resetn, stream_source_dpi_bfm_relu1_out0_inst:resetn, stream_source_dpi_bfm_relu2_in0_inst:resetn, stream_source_dpi_bfm_relu2_out0_inst:resetn, stream_source_dpi_bfm_relu3_in0_inst:resetn, stream_source_dpi_bfm_relu3_out0_inst:resetn, stream_source_dpi_bfm_relu4_in0_inst:resetn, stream_source_dpi_bfm_relu4_out0_inst:resetn, stream_source_dpi_bfm_softmax_in0_inst:resetn, stream_source_dpi_bfm_softmax_out0_inst:resetn]
	wire         component_dpi_controller_avgpooling1_inst_component_irq_irq;                                   // irq_mapper:sender_irq -> component_dpi_controller_avgpooling1_inst:done_irq
	wire         component_dpi_controller_avgpooling2_inst_component_irq_irq;                                   // irq_mapper_001:sender_irq -> component_dpi_controller_avgpooling2_inst:done_irq
	wire         component_dpi_controller_conv1_inst_component_irq_irq;                                         // irq_mapper_002:sender_irq -> component_dpi_controller_conv1_inst:done_irq
	wire         component_dpi_controller_conv2_inst_component_irq_irq;                                         // irq_mapper_003:sender_irq -> component_dpi_controller_conv2_inst:done_irq
	wire         component_dpi_controller_fc1_inst_component_irq_irq;                                           // irq_mapper_004:sender_irq -> component_dpi_controller_fc1_inst:done_irq
	wire         component_dpi_controller_fc3_inst_component_irq_irq;                                           // irq_mapper_005:sender_irq -> component_dpi_controller_fc3_inst:done_irq
	wire         component_dpi_controller_relu1_inst_component_irq_irq;                                         // irq_mapper_006:sender_irq -> component_dpi_controller_relu1_inst:done_irq
	wire         component_dpi_controller_relu2_inst_component_irq_irq;                                         // irq_mapper_007:sender_irq -> component_dpi_controller_relu2_inst:done_irq
	wire         component_dpi_controller_relu3_inst_component_irq_irq;                                         // irq_mapper_008:sender_irq -> component_dpi_controller_relu3_inst:done_irq
	wire         component_dpi_controller_relu4_inst_component_irq_irq;                                         // irq_mapper_009:sender_irq -> component_dpi_controller_relu4_inst:done_irq
	wire         component_dpi_controller_softmax_inst_component_irq_irq;                                       // irq_mapper_010:sender_irq -> component_dpi_controller_softmax_inst:done_irq

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst avgpooling1_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_avgpooling1_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (avgpooling1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (avgpooling1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (avgpooling1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst avgpooling1_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_avgpooling1_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (avgpooling1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (avgpooling1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (avgpooling1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_avgpooling1_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit)  // out_conduit_1.conduit
	);

	tb_avgpooling1_inst avgpooling1_inst (
		.avmm_0_rw_address    (avgpooling1_inst_avmm_0_rw_address),                               // avmm_0_rw.address
		.avmm_0_rw_byteenable (avgpooling1_inst_avmm_0_rw_byteenable),                            //          .byteenable
		.avmm_0_rw_read       (avgpooling1_inst_avmm_0_rw_read),                                  //          .read
		.avmm_0_rw_readdata   (avgpooling1_inst_avmm_0_rw_readdata),                              //          .readdata
		.avmm_0_rw_write      (avgpooling1_inst_avmm_0_rw_write),                                 //          .write
		.avmm_0_rw_writedata  (avgpooling1_inst_avmm_0_rw_writedata),                             //          .writedata
		.start                (component_dpi_controller_avgpooling1_inst_component_call_valid),   //      call.valid
		.busy                 (avgpooling1_inst_call_stall),                                      //          .stall
		.clock                (clock_reset_inst_clock_clk),                                       //     clock.clk
		.in0                  (stream_source_dpi_bfm_avgpooling1_in0_inst_source_data_data),      //       in0.data
		.out0                 (stream_source_dpi_bfm_avgpooling1_out0_inst_source_data_data),     //      out0.data
		.resetn               (clock_reset_inst_reset_reset),                                     //     reset.reset_n
		.done                 (avgpooling1_inst_return_valid),                                    //    return.valid
		.stall                (component_dpi_controller_avgpooling1_inst_component_return_stall)  //          .stall
	);

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst avgpooling2_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_avgpooling2_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (avgpooling2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (avgpooling2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (avgpooling2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst avgpooling2_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_avgpooling2_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (avgpooling2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (avgpooling2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (avgpooling2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst avgpooling2_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_avgpooling2_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (avgpooling2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (avgpooling2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit)  // out_conduit_1.conduit
	);

	tb_avgpooling2_inst avgpooling2_inst (
		.avmm_0_rw_address    (avgpooling2_inst_avmm_0_rw_address),                               // avmm_0_rw.address
		.avmm_0_rw_byteenable (avgpooling2_inst_avmm_0_rw_byteenable),                            //          .byteenable
		.avmm_0_rw_read       (avgpooling2_inst_avmm_0_rw_read),                                  //          .read
		.avmm_0_rw_readdata   (avgpooling2_inst_avmm_0_rw_readdata),                              //          .readdata
		.avmm_0_rw_write      (avgpooling2_inst_avmm_0_rw_write),                                 //          .write
		.avmm_0_rw_writedata  (avgpooling2_inst_avmm_0_rw_writedata),                             //          .writedata
		.start                (component_dpi_controller_avgpooling2_inst_component_call_valid),   //      call.valid
		.busy                 (avgpooling2_inst_call_stall),                                      //          .stall
		.clock                (clock_reset_inst_clock_clk),                                       //     clock.clk
		.in0                  (stream_source_dpi_bfm_avgpooling2_in0_inst_source_data_data),      //       in0.data
		.out0                 (stream_source_dpi_bfm_avgpooling2_out0_inst_source_data_data),     //      out0.data
		.resetn               (clock_reset_inst_reset_reset),                                     //     reset.reset_n
		.done                 (avgpooling2_inst_return_valid),                                    //    return.valid
		.stall                (component_dpi_controller_avgpooling2_inst_component_return_stall)  //          .stall
	);

	hls_sim_clock_reset #(
		.RESET_CYCLE_HOLD (4)
	) clock_reset_inst (
		.clock         (clock_reset_inst_clock_clk),                  //      clock.clk
		.resetn        (clock_reset_inst_reset_reset),                //      reset.reset_n
		.clock2x       (clock_reset_inst_clock2x_clk),                //    clock2x.clk
		.trigger_reset (main_dpi_controller_inst_reset_ctrl_conduit)  // reset_ctrl.conduit
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("avgpooling1"),
		.COMPONENT_MANGLED_NAME       ("\\3favgpooling1@@YAXQEAY1BM@BM@MQEAY1O@O@M@Z"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_avgpooling1_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                         //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                       //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                       //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_avgpooling1_inst_dpi_control_bind_conduit),                 //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_avgpooling1_inst_dpi_control_enable_conduit),               //               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_0_conduit),                                   //                component_enabled.conduit
		.component_done                   (component_dpi_controller_avgpooling1_inst_component_done_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_avgpooling1_inst_component_wait_for_stream_writes_conduit), // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                                   //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_avgpooling1_inst_read_implicit_streams_conduit),            //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                                   //             readback_from_agents.conduit
		.start                            (component_dpi_controller_avgpooling1_inst_component_call_valid),                     //                   component_call.valid
		.busy                             (avgpooling1_inst_call_stall),                                                        //                                 .stall
		.done                             (avgpooling1_inst_return_valid),                                                      //                 component_return.valid
		.stall                            (component_dpi_controller_avgpooling1_inst_component_return_stall),                   //                                 .stall
		.done_irq                         (component_dpi_controller_avgpooling1_inst_component_irq_irq),                        //                    component_irq.irq
		.returndata                       ()                                                                                    //                       returndata.data
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("avgpooling2"),
		.COMPONENT_MANGLED_NAME       ("\\3favgpooling2@@YAXQEAY199MQEAY144M@Z"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_avgpooling2_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                         //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                       //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                       //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_avgpooling2_inst_dpi_control_bind_conduit),                 //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_avgpooling2_inst_dpi_control_enable_conduit),               //               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_1_conduit),                                   //                component_enabled.conduit
		.component_done                   (component_dpi_controller_avgpooling2_inst_component_done_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_avgpooling2_inst_component_wait_for_stream_writes_conduit), // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                                   //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_avgpooling2_inst_read_implicit_streams_conduit),            //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                                   //             readback_from_agents.conduit
		.start                            (component_dpi_controller_avgpooling2_inst_component_call_valid),                     //                   component_call.valid
		.busy                             (avgpooling2_inst_call_stall),                                                        //                                 .stall
		.done                             (avgpooling2_inst_return_valid),                                                      //                 component_return.valid
		.stall                            (component_dpi_controller_avgpooling2_inst_component_return_stall),                   //                                 .stall
		.done_irq                         (component_dpi_controller_avgpooling2_inst_component_irq_irq),                        //                    component_irq.irq
		.returndata                       ()                                                                                    //                       returndata.data
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("conv1"),
		.COMPONENT_MANGLED_NAME       ("\\3fconv1@@YAXQEAY0BM@MQEAY100MQEAMQEAY1BM@BM@M@Z"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_conv1_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                   //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                 //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                 //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_conv1_inst_dpi_control_bind_conduit),                 //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_conv1_inst_dpi_control_enable_conduit),               //               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_2_conduit),                             //                component_enabled.conduit
		.component_done                   (component_dpi_controller_conv1_inst_component_done_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_conv1_inst_component_wait_for_stream_writes_conduit), // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                             //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_conv1_inst_read_implicit_streams_conduit),            //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                             //             readback_from_agents.conduit
		.start                            (component_dpi_controller_conv1_inst_component_call_valid),                     //                   component_call.valid
		.busy                             (conv1_inst_call_stall),                                                        //                                 .stall
		.done                             (conv1_inst_return_valid),                                                      //                 component_return.valid
		.stall                            (component_dpi_controller_conv1_inst_component_return_stall),                   //                                 .stall
		.done_irq                         (component_dpi_controller_conv1_inst_component_irq_irq),                        //                    component_irq.irq
		.returndata                       ()                                                                              //                       returndata.data
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("conv2"),
		.COMPONENT_MANGLED_NAME       ("\\3fconv2@@YAXQEAY1O@O@MQEAY2544MQEAMQEAY199M@Z"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_conv2_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                   //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                 //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                 //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_conv2_inst_dpi_control_bind_conduit),                 //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_conv2_inst_dpi_control_enable_conduit),               //               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_3_conduit),                             //                component_enabled.conduit
		.component_done                   (component_dpi_controller_conv2_inst_component_done_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_conv2_inst_component_wait_for_stream_writes_conduit), // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                             //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_conv2_inst_read_implicit_streams_conduit),            //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                             //             readback_from_agents.conduit
		.start                            (component_dpi_controller_conv2_inst_component_call_valid),                     //                   component_call.valid
		.busy                             (conv2_inst_call_stall),                                                        //                                 .stall
		.done                             (conv2_inst_return_valid),                                                      //                 component_return.valid
		.stall                            (component_dpi_controller_conv2_inst_component_return_stall),                   //                                 .stall
		.done_irq                         (component_dpi_controller_conv2_inst_component_irq_irq),                        //                    component_irq.irq
		.returndata                       ()                                                                              //                       returndata.data
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("fc1"),
		.COMPONENT_MANGLED_NAME       ("\\3ffc1@@YAXQEAMQEAY0BJA@M00@Z"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_fc1_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                 //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                               //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                               //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_fc1_inst_dpi_control_bind_conduit),                 //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_fc1_inst_dpi_control_enable_conduit),               //               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_4_conduit),                           //                component_enabled.conduit
		.component_done                   (component_dpi_controller_fc1_inst_component_done_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_fc1_inst_component_wait_for_stream_writes_conduit), // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                           //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_fc1_inst_read_implicit_streams_conduit),            //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                           //             readback_from_agents.conduit
		.start                            (component_dpi_controller_fc1_inst_component_call_valid),                     //                   component_call.valid
		.busy                             (fc1_inst_call_stall),                                                        //                                 .stall
		.done                             (fc1_inst_return_valid),                                                      //                 component_return.valid
		.stall                            (component_dpi_controller_fc1_inst_component_return_stall),                   //                                 .stall
		.done_irq                         (component_dpi_controller_fc1_inst_component_irq_irq),                        //                    component_irq.irq
		.returndata                       ()                                                                            //                       returndata.data
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("fc3"),
		.COMPONENT_MANGLED_NAME       ("\\3ffc3@@YAXQEAMQEAY0FE@M00@Z"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_fc3_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                 //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                               //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                               //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_fc3_inst_dpi_control_bind_conduit),                 //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_fc3_inst_dpi_control_enable_conduit),               //               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_5_conduit),                           //                component_enabled.conduit
		.component_done                   (component_dpi_controller_fc3_inst_component_done_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_fc3_inst_component_wait_for_stream_writes_conduit), // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                           //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_fc3_inst_read_implicit_streams_conduit),            //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                           //             readback_from_agents.conduit
		.start                            (component_dpi_controller_fc3_inst_component_call_valid),                     //                   component_call.valid
		.busy                             (fc3_inst_call_stall),                                                        //                                 .stall
		.done                             (fc3_inst_return_valid),                                                      //                 component_return.valid
		.stall                            (component_dpi_controller_fc3_inst_component_return_stall),                   //                                 .stall
		.done_irq                         (component_dpi_controller_fc3_inst_component_irq_irq),                        //                    component_irq.irq
		.returndata                       ()                                                                            //                       returndata.data
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("relu1"),
		.COMPONENT_MANGLED_NAME       ("\\3frelu1@@YAXQEAY1BM@BM@M0@Z"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_relu1_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                   //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                 //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                 //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_relu1_inst_dpi_control_bind_conduit),                 //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_relu1_inst_dpi_control_enable_conduit),               //               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_6_conduit),                             //                component_enabled.conduit
		.component_done                   (component_dpi_controller_relu1_inst_component_done_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_relu1_inst_component_wait_for_stream_writes_conduit), // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                             //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_relu1_inst_read_implicit_streams_conduit),            //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                             //             readback_from_agents.conduit
		.start                            (component_dpi_controller_relu1_inst_component_call_valid),                     //                   component_call.valid
		.busy                             (relu1_inst_call_stall),                                                        //                                 .stall
		.done                             (relu1_inst_return_valid),                                                      //                 component_return.valid
		.stall                            (component_dpi_controller_relu1_inst_component_return_stall),                   //                                 .stall
		.done_irq                         (component_dpi_controller_relu1_inst_component_irq_irq),                        //                    component_irq.irq
		.returndata                       ()                                                                              //                       returndata.data
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("relu2"),
		.COMPONENT_MANGLED_NAME       ("\\3frelu2@@YAXQEAY199M0@Z"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_relu2_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                   //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                 //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                 //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_relu2_inst_dpi_control_bind_conduit),                 //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_relu2_inst_dpi_control_enable_conduit),               //               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_7_conduit),                             //                component_enabled.conduit
		.component_done                   (component_dpi_controller_relu2_inst_component_done_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_relu2_inst_component_wait_for_stream_writes_conduit), // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                             //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_relu2_inst_read_implicit_streams_conduit),            //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                             //             readback_from_agents.conduit
		.start                            (component_dpi_controller_relu2_inst_component_call_valid),                     //                   component_call.valid
		.busy                             (relu2_inst_call_stall),                                                        //                                 .stall
		.done                             (relu2_inst_return_valid),                                                      //                 component_return.valid
		.stall                            (component_dpi_controller_relu2_inst_component_return_stall),                   //                                 .stall
		.done_irq                         (component_dpi_controller_relu2_inst_component_irq_irq),                        //                    component_irq.irq
		.returndata                       ()                                                                              //                       returndata.data
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("relu3"),
		.COMPONENT_MANGLED_NAME       ("\\3frelu3@@YAXQEAM0@Z"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_relu3_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                   //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                 //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                 //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_relu3_inst_dpi_control_bind_conduit),                 //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_relu3_inst_dpi_control_enable_conduit),               //               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_8_conduit),                             //                component_enabled.conduit
		.component_done                   (component_dpi_controller_relu3_inst_component_done_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_relu3_inst_component_wait_for_stream_writes_conduit), // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                             //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_relu3_inst_read_implicit_streams_conduit),            //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                             //             readback_from_agents.conduit
		.start                            (component_dpi_controller_relu3_inst_component_call_valid),                     //                   component_call.valid
		.busy                             (relu3_inst_call_stall),                                                        //                                 .stall
		.done                             (relu3_inst_return_valid),                                                      //                 component_return.valid
		.stall                            (component_dpi_controller_relu3_inst_component_return_stall),                   //                                 .stall
		.done_irq                         (component_dpi_controller_relu3_inst_component_irq_irq),                        //                    component_irq.irq
		.returndata                       ()                                                                              //                       returndata.data
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("relu4"),
		.COMPONENT_MANGLED_NAME       ("\\3frelu4@@YAXQEAM0@Z"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_relu4_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                   //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                 //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                 //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_relu4_inst_dpi_control_bind_conduit),                 //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_relu4_inst_dpi_control_enable_conduit),               //               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_9_conduit),                             //                component_enabled.conduit
		.component_done                   (component_dpi_controller_relu4_inst_component_done_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_relu4_inst_component_wait_for_stream_writes_conduit), // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                             //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_relu4_inst_read_implicit_streams_conduit),            //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                             //             readback_from_agents.conduit
		.start                            (component_dpi_controller_relu4_inst_component_call_valid),                     //                   component_call.valid
		.busy                             (relu4_inst_call_stall),                                                        //                                 .stall
		.done                             (relu4_inst_return_valid),                                                      //                 component_return.valid
		.stall                            (component_dpi_controller_relu4_inst_component_return_stall),                   //                                 .stall
		.done_irq                         (component_dpi_controller_relu4_inst_component_irq_irq),                        //                    component_irq.irq
		.returndata                       ()                                                                              //                       returndata.data
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("softmax"),
		.COMPONENT_MANGLED_NAME       ("\\3fsoftmax@@YAXQEAM0@Z"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_softmax_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                     //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                   //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                   //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_softmax_inst_dpi_control_bind_conduit),                 //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_softmax_inst_dpi_control_enable_conduit),               //               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_10_conduit),                              //                component_enabled.conduit
		.component_done                   (component_dpi_controller_softmax_inst_component_done_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_softmax_inst_component_wait_for_stream_writes_conduit), // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                               //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_softmax_inst_read_implicit_streams_conduit),            //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                               //             readback_from_agents.conduit
		.start                            (component_dpi_controller_softmax_inst_component_call_valid),                     //                   component_call.valid
		.busy                             (softmax_inst_call_stall),                                                        //                                 .stall
		.done                             (softmax_inst_return_valid),                                                      //                 component_return.valid
		.stall                            (component_dpi_controller_softmax_inst_component_return_stall),                   //                                 .stall
		.done_irq                         (component_dpi_controller_softmax_inst_component_irq_irq),                        //                    component_irq.irq
		.returndata                       ()                                                                                //                       returndata.data
	);

	tb_concatenate_component_done_inst concatenate_component_done_inst (
		.out_conduit   (concatenate_component_done_inst_out_conduit_conduit),              //   out_conduit.conduit
		.in_conduit_0  (component_dpi_controller_avgpooling1_inst_component_done_conduit), //  in_conduit_0.conduit
		.in_conduit_1  (component_dpi_controller_avgpooling2_inst_component_done_conduit), //  in_conduit_1.conduit
		.in_conduit_2  (component_dpi_controller_conv1_inst_component_done_conduit),       //  in_conduit_2.conduit
		.in_conduit_3  (component_dpi_controller_conv2_inst_component_done_conduit),       //  in_conduit_3.conduit
		.in_conduit_4  (component_dpi_controller_fc1_inst_component_done_conduit),         //  in_conduit_4.conduit
		.in_conduit_5  (component_dpi_controller_fc3_inst_component_done_conduit),         //  in_conduit_5.conduit
		.in_conduit_6  (component_dpi_controller_relu1_inst_component_done_conduit),       //  in_conduit_6.conduit
		.in_conduit_7  (component_dpi_controller_relu2_inst_component_done_conduit),       //  in_conduit_7.conduit
		.in_conduit_8  (component_dpi_controller_relu3_inst_component_done_conduit),       //  in_conduit_8.conduit
		.in_conduit_9  (component_dpi_controller_relu4_inst_component_done_conduit),       //  in_conduit_9.conduit
		.in_conduit_10 (component_dpi_controller_softmax_inst_component_done_conduit)      // in_conduit_10.conduit
	);

	tb_concatenate_component_done_inst concatenate_component_wait_for_stream_writes_inst (
		.out_conduit   (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit),              //   out_conduit.conduit
		.in_conduit_0  (component_dpi_controller_avgpooling1_inst_component_wait_for_stream_writes_conduit), //  in_conduit_0.conduit
		.in_conduit_1  (component_dpi_controller_avgpooling2_inst_component_wait_for_stream_writes_conduit), //  in_conduit_1.conduit
		.in_conduit_2  (component_dpi_controller_conv1_inst_component_wait_for_stream_writes_conduit),       //  in_conduit_2.conduit
		.in_conduit_3  (component_dpi_controller_conv2_inst_component_wait_for_stream_writes_conduit),       //  in_conduit_3.conduit
		.in_conduit_4  (component_dpi_controller_fc1_inst_component_wait_for_stream_writes_conduit),         //  in_conduit_4.conduit
		.in_conduit_5  (component_dpi_controller_fc3_inst_component_wait_for_stream_writes_conduit),         //  in_conduit_5.conduit
		.in_conduit_6  (component_dpi_controller_relu1_inst_component_wait_for_stream_writes_conduit),       //  in_conduit_6.conduit
		.in_conduit_7  (component_dpi_controller_relu2_inst_component_wait_for_stream_writes_conduit),       //  in_conduit_7.conduit
		.in_conduit_8  (component_dpi_controller_relu3_inst_component_wait_for_stream_writes_conduit),       //  in_conduit_8.conduit
		.in_conduit_9  (component_dpi_controller_relu4_inst_component_wait_for_stream_writes_conduit),       //  in_conduit_9.conduit
		.in_conduit_10 (component_dpi_controller_softmax_inst_component_wait_for_stream_writes_conduit)      // in_conduit_10.conduit
	);

	tb_conv1_component_dpi_controller_bind_conduit_fanout_inst conv1_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_conv1_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit), // out_conduit_3.conduit
		.out_conduit_4 (conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit)  // out_conduit_4.conduit
	);

	tb_conv1_component_dpi_controller_bind_conduit_fanout_inst conv1_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_conv1_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit), // out_conduit_3.conduit
		.out_conduit_4 (conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit)  // out_conduit_4.conduit
	);

	tb_conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_conv1_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit)  // out_conduit_3.conduit
	);

	tb_conv1_inst conv1_inst (
		.avmm_0_rw_address    (conv1_inst_avmm_0_rw_address),                               // avmm_0_rw.address
		.avmm_0_rw_byteenable (conv1_inst_avmm_0_rw_byteenable),                            //          .byteenable
		.avmm_0_rw_read       (conv1_inst_avmm_0_rw_read),                                  //          .read
		.avmm_0_rw_readdata   (conv1_inst_avmm_0_rw_readdata),                              //          .readdata
		.avmm_0_rw_write      (conv1_inst_avmm_0_rw_write),                                 //          .write
		.avmm_0_rw_writedata  (conv1_inst_avmm_0_rw_writedata),                             //          .writedata
		.bias                 (stream_source_dpi_bfm_conv1_bias_inst_source_data_data),     //      bias.data
		.start                (component_dpi_controller_conv1_inst_component_call_valid),   //      call.valid
		.busy                 (conv1_inst_call_stall),                                      //          .stall
		.clock                (clock_reset_inst_clock_clk),                                 //     clock.clk
		.in0                  (stream_source_dpi_bfm_conv1_in0_inst_source_data_data),      //       in0.data
		.kernel               (stream_source_dpi_bfm_conv1_kernel_inst_source_data_data),   //    kernel.data
		.out0                 (stream_source_dpi_bfm_conv1_out0_inst_source_data_data),     //      out0.data
		.resetn               (clock_reset_inst_reset_reset),                               //     reset.reset_n
		.done                 (conv1_inst_return_valid),                                    //    return.valid
		.stall                (component_dpi_controller_conv1_inst_component_return_stall)  //          .stall
	);

	tb_conv1_component_dpi_controller_bind_conduit_fanout_inst conv2_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_conv2_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit), // out_conduit_3.conduit
		.out_conduit_4 (conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit)  // out_conduit_4.conduit
	);

	tb_conv1_component_dpi_controller_bind_conduit_fanout_inst conv2_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_conv2_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit), // out_conduit_3.conduit
		.out_conduit_4 (conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit)  // out_conduit_4.conduit
	);

	tb_conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_conv2_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit)  // out_conduit_3.conduit
	);

	tb_conv2_inst conv2_inst (
		.avmm_0_rw_address    (conv2_inst_avmm_0_rw_address),                               // avmm_0_rw.address
		.avmm_0_rw_byteenable (conv2_inst_avmm_0_rw_byteenable),                            //          .byteenable
		.avmm_0_rw_read       (conv2_inst_avmm_0_rw_read),                                  //          .read
		.avmm_0_rw_readdata   (conv2_inst_avmm_0_rw_readdata),                              //          .readdata
		.avmm_0_rw_write      (conv2_inst_avmm_0_rw_write),                                 //          .write
		.avmm_0_rw_writedata  (conv2_inst_avmm_0_rw_writedata),                             //          .writedata
		.bias                 (stream_source_dpi_bfm_conv2_bias_inst_source_data_data),     //      bias.data
		.start                (component_dpi_controller_conv2_inst_component_call_valid),   //      call.valid
		.busy                 (conv2_inst_call_stall),                                      //          .stall
		.clock                (clock_reset_inst_clock_clk),                                 //     clock.clk
		.in0                  (stream_source_dpi_bfm_conv2_in0_inst_source_data_data),      //       in0.data
		.kernel               (stream_source_dpi_bfm_conv2_kernel_inst_source_data_data),   //    kernel.data
		.out0                 (stream_source_dpi_bfm_conv2_out0_inst_source_data_data),     //      out0.data
		.resetn               (clock_reset_inst_reset_reset),                               //     reset.reset_n
		.done                 (conv2_inst_return_valid),                                    //    return.valid
		.stall                (component_dpi_controller_conv2_inst_component_return_stall)  //          .stall
	);

	tb_conv1_component_dpi_controller_bind_conduit_fanout_inst fc1_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_fc1_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit), // out_conduit_3.conduit
		.out_conduit_4 (fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit)  // out_conduit_4.conduit
	);

	tb_conv1_component_dpi_controller_bind_conduit_fanout_inst fc1_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_fc1_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit), // out_conduit_3.conduit
		.out_conduit_4 (fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit)  // out_conduit_4.conduit
	);

	tb_conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_fc1_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit)  // out_conduit_3.conduit
	);

	tb_fc1_inst fc1_inst (
		.avmm_0_rw_address    (fc1_inst_avmm_0_rw_address),                               // avmm_0_rw.address
		.avmm_0_rw_byteenable (fc1_inst_avmm_0_rw_byteenable),                            //          .byteenable
		.avmm_0_rw_read       (fc1_inst_avmm_0_rw_read),                                  //          .read
		.avmm_0_rw_readdata   (fc1_inst_avmm_0_rw_readdata),                              //          .readdata
		.avmm_0_rw_write      (fc1_inst_avmm_0_rw_write),                                 //          .write
		.avmm_0_rw_writedata  (fc1_inst_avmm_0_rw_writedata),                             //          .writedata
		.bias                 (stream_source_dpi_bfm_fc1_bias_inst_source_data_data),     //      bias.data
		.start                (component_dpi_controller_fc1_inst_component_call_valid),   //      call.valid
		.busy                 (fc1_inst_call_stall),                                      //          .stall
		.clock                (clock_reset_inst_clock_clk),                               //     clock.clk
		.in0                  (stream_source_dpi_bfm_fc1_in0_inst_source_data_data),      //       in0.data
		.out0                 (stream_source_dpi_bfm_fc1_out0_inst_source_data_data),     //      out0.data
		.resetn               (clock_reset_inst_reset_reset),                             //     reset.reset_n
		.done                 (fc1_inst_return_valid),                                    //    return.valid
		.stall                (component_dpi_controller_fc1_inst_component_return_stall), //          .stall
		.weights              (stream_source_dpi_bfm_fc1_weights_inst_source_data_data)   //   weights.data
	);

	tb_conv1_component_dpi_controller_bind_conduit_fanout_inst fc3_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_fc3_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit), // out_conduit_3.conduit
		.out_conduit_4 (fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit)  // out_conduit_4.conduit
	);

	tb_conv1_component_dpi_controller_bind_conduit_fanout_inst fc3_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_fc3_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit), // out_conduit_3.conduit
		.out_conduit_4 (fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit)  // out_conduit_4.conduit
	);

	tb_conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_fc3_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit)  // out_conduit_3.conduit
	);

	tb_fc3_inst fc3_inst (
		.avmm_0_rw_address    (fc3_inst_avmm_0_rw_address),                               // avmm_0_rw.address
		.avmm_0_rw_byteenable (fc3_inst_avmm_0_rw_byteenable),                            //          .byteenable
		.avmm_0_rw_read       (fc3_inst_avmm_0_rw_read),                                  //          .read
		.avmm_0_rw_readdata   (fc3_inst_avmm_0_rw_readdata),                              //          .readdata
		.avmm_0_rw_write      (fc3_inst_avmm_0_rw_write),                                 //          .write
		.avmm_0_rw_writedata  (fc3_inst_avmm_0_rw_writedata),                             //          .writedata
		.bias                 (stream_source_dpi_bfm_fc3_bias_inst_source_data_data),     //      bias.data
		.start                (component_dpi_controller_fc3_inst_component_call_valid),   //      call.valid
		.busy                 (fc3_inst_call_stall),                                      //          .stall
		.clock                (clock_reset_inst_clock_clk),                               //     clock.clk
		.in0                  (stream_source_dpi_bfm_fc3_in0_inst_source_data_data),      //       in0.data
		.out0                 (stream_source_dpi_bfm_fc3_out0_inst_source_data_data),     //      out0.data
		.resetn               (clock_reset_inst_reset_reset),                             //     reset.reset_n
		.done                 (fc3_inst_return_valid),                                    //    return.valid
		.stall                (component_dpi_controller_fc3_inst_component_return_stall), //          .stall
		.weights              (stream_source_dpi_bfm_fc3_weights_inst_source_data_data)   //   weights.data
	);

	hls_sim_main_dpi_controller #(
		.NUM_COMPONENTS      (11),
		.COMPONENT_NAMES_STR ("avgpooling1,avgpooling2,conv1,conv2,fc1,fc3,relu1,relu2,relu3,relu4,softmax")
	) main_dpi_controller_inst (
		.clock                            (clock_reset_inst_clock_clk),                                            //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                          //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                          //                          clock2x.clk
		.component_enabled                (main_dpi_controller_inst_component_enabled_conduit),                    //                component_enabled.conduit
		.component_done                   (concatenate_component_done_inst_out_conduit_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit), // component_wait_for_stream_writes.conduit
		.trigger_reset                    (main_dpi_controller_inst_reset_ctrl_conduit)                            //                       reset_ctrl.conduit
	);

	hls_sim_mm_agent_dpi_bfm #(
		.AV_ADDRESS_W               (64),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (8),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.COMPONENT_NAME             ("avgpooling1"),
		.INTERFACE_ID               (0)
	) mm_agent_dpi_bfm_avgpooling1_avmm_0_rw_inst (
		.do_bind           (avgpooling1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),   //   dpi_control_bind.conduit
		.enable            (avgpooling1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // dpi_control_enable.conduit
		.clock             (clock_reset_inst_clock_clk),                                                            //              clock.clk
		.reset_n           (clock_reset_inst_reset_reset),                                                          //              reset.reset_n
		.avs_writedata     (avgpooling1_inst_avmm_0_rw_writedata),                                                  //                 s0.writedata
		.avs_readdata      (avgpooling1_inst_avmm_0_rw_readdata),                                                   //                   .readdata
		.avs_address       (avgpooling1_inst_avmm_0_rw_address),                                                    //                   .address
		.avs_write         (avgpooling1_inst_avmm_0_rw_write),                                                      //                   .write
		.avs_read          (avgpooling1_inst_avmm_0_rw_read),                                                       //                   .read
		.avs_byteenable    (avgpooling1_inst_avmm_0_rw_byteenable),                                                 //                   .byteenable
		.avs_readdatavalid ()                                                                                       //        (terminated)
	);

	hls_sim_mm_agent_dpi_bfm #(
		.AV_ADDRESS_W               (64),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (8),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.COMPONENT_NAME             ("avgpooling2"),
		.INTERFACE_ID               (0)
	) mm_agent_dpi_bfm_avgpooling2_avmm_0_rw_inst (
		.do_bind           (avgpooling2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),   //   dpi_control_bind.conduit
		.enable            (avgpooling2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // dpi_control_enable.conduit
		.clock             (clock_reset_inst_clock_clk),                                                            //              clock.clk
		.reset_n           (clock_reset_inst_reset_reset),                                                          //              reset.reset_n
		.avs_writedata     (avgpooling2_inst_avmm_0_rw_writedata),                                                  //                 s0.writedata
		.avs_readdata      (avgpooling2_inst_avmm_0_rw_readdata),                                                   //                   .readdata
		.avs_address       (avgpooling2_inst_avmm_0_rw_address),                                                    //                   .address
		.avs_write         (avgpooling2_inst_avmm_0_rw_write),                                                      //                   .write
		.avs_read          (avgpooling2_inst_avmm_0_rw_read),                                                       //                   .read
		.avs_byteenable    (avgpooling2_inst_avmm_0_rw_byteenable),                                                 //                   .byteenable
		.avs_readdatavalid ()                                                                                       //        (terminated)
	);

	hls_sim_mm_agent_dpi_bfm #(
		.AV_ADDRESS_W               (64),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (8),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.COMPONENT_NAME             ("conv1"),
		.INTERFACE_ID               (0)
	) mm_agent_dpi_bfm_conv1_avmm_0_rw_inst (
		.do_bind           (conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),   //   dpi_control_bind.conduit
		.enable            (conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // dpi_control_enable.conduit
		.clock             (clock_reset_inst_clock_clk),                                                      //              clock.clk
		.reset_n           (clock_reset_inst_reset_reset),                                                    //              reset.reset_n
		.avs_writedata     (conv1_inst_avmm_0_rw_writedata),                                                  //                 s0.writedata
		.avs_readdata      (conv1_inst_avmm_0_rw_readdata),                                                   //                   .readdata
		.avs_address       (conv1_inst_avmm_0_rw_address),                                                    //                   .address
		.avs_write         (conv1_inst_avmm_0_rw_write),                                                      //                   .write
		.avs_read          (conv1_inst_avmm_0_rw_read),                                                       //                   .read
		.avs_byteenable    (conv1_inst_avmm_0_rw_byteenable),                                                 //                   .byteenable
		.avs_readdatavalid ()                                                                                 //        (terminated)
	);

	hls_sim_mm_agent_dpi_bfm #(
		.AV_ADDRESS_W               (64),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (8),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.COMPONENT_NAME             ("conv2"),
		.INTERFACE_ID               (0)
	) mm_agent_dpi_bfm_conv2_avmm_0_rw_inst (
		.do_bind           (conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),   //   dpi_control_bind.conduit
		.enable            (conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // dpi_control_enable.conduit
		.clock             (clock_reset_inst_clock_clk),                                                      //              clock.clk
		.reset_n           (clock_reset_inst_reset_reset),                                                    //              reset.reset_n
		.avs_writedata     (conv2_inst_avmm_0_rw_writedata),                                                  //                 s0.writedata
		.avs_readdata      (conv2_inst_avmm_0_rw_readdata),                                                   //                   .readdata
		.avs_address       (conv2_inst_avmm_0_rw_address),                                                    //                   .address
		.avs_write         (conv2_inst_avmm_0_rw_write),                                                      //                   .write
		.avs_read          (conv2_inst_avmm_0_rw_read),                                                       //                   .read
		.avs_byteenable    (conv2_inst_avmm_0_rw_byteenable),                                                 //                   .byteenable
		.avs_readdatavalid ()                                                                                 //        (terminated)
	);

	hls_sim_mm_agent_dpi_bfm #(
		.AV_ADDRESS_W               (64),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (8),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.COMPONENT_NAME             ("fc1"),
		.INTERFACE_ID               (0)
	) mm_agent_dpi_bfm_fc1_avmm_0_rw_inst (
		.do_bind           (fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),   //   dpi_control_bind.conduit
		.enable            (fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // dpi_control_enable.conduit
		.clock             (clock_reset_inst_clock_clk),                                                    //              clock.clk
		.reset_n           (clock_reset_inst_reset_reset),                                                  //              reset.reset_n
		.avs_writedata     (fc1_inst_avmm_0_rw_writedata),                                                  //                 s0.writedata
		.avs_readdata      (fc1_inst_avmm_0_rw_readdata),                                                   //                   .readdata
		.avs_address       (fc1_inst_avmm_0_rw_address),                                                    //                   .address
		.avs_write         (fc1_inst_avmm_0_rw_write),                                                      //                   .write
		.avs_read          (fc1_inst_avmm_0_rw_read),                                                       //                   .read
		.avs_byteenable    (fc1_inst_avmm_0_rw_byteenable),                                                 //                   .byteenable
		.avs_readdatavalid ()                                                                               //        (terminated)
	);

	hls_sim_mm_agent_dpi_bfm #(
		.AV_ADDRESS_W               (64),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (8),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.COMPONENT_NAME             ("fc3"),
		.INTERFACE_ID               (0)
	) mm_agent_dpi_bfm_fc3_avmm_0_rw_inst (
		.do_bind           (fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),   //   dpi_control_bind.conduit
		.enable            (fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // dpi_control_enable.conduit
		.clock             (clock_reset_inst_clock_clk),                                                    //              clock.clk
		.reset_n           (clock_reset_inst_reset_reset),                                                  //              reset.reset_n
		.avs_writedata     (fc3_inst_avmm_0_rw_writedata),                                                  //                 s0.writedata
		.avs_readdata      (fc3_inst_avmm_0_rw_readdata),                                                   //                   .readdata
		.avs_address       (fc3_inst_avmm_0_rw_address),                                                    //                   .address
		.avs_write         (fc3_inst_avmm_0_rw_write),                                                      //                   .write
		.avs_read          (fc3_inst_avmm_0_rw_read),                                                       //                   .read
		.avs_byteenable    (fc3_inst_avmm_0_rw_byteenable),                                                 //                   .byteenable
		.avs_readdatavalid ()                                                                               //        (terminated)
	);

	hls_sim_mm_agent_dpi_bfm #(
		.AV_ADDRESS_W               (64),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (8),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.COMPONENT_NAME             ("relu1"),
		.INTERFACE_ID               (0)
	) mm_agent_dpi_bfm_relu1_avmm_0_rw_inst (
		.do_bind           (relu1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),   //   dpi_control_bind.conduit
		.enable            (relu1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // dpi_control_enable.conduit
		.clock             (clock_reset_inst_clock_clk),                                                      //              clock.clk
		.reset_n           (clock_reset_inst_reset_reset),                                                    //              reset.reset_n
		.avs_writedata     (relu1_inst_avmm_0_rw_writedata),                                                  //                 s0.writedata
		.avs_readdata      (relu1_inst_avmm_0_rw_readdata),                                                   //                   .readdata
		.avs_address       (relu1_inst_avmm_0_rw_address),                                                    //                   .address
		.avs_write         (relu1_inst_avmm_0_rw_write),                                                      //                   .write
		.avs_read          (relu1_inst_avmm_0_rw_read),                                                       //                   .read
		.avs_byteenable    (relu1_inst_avmm_0_rw_byteenable),                                                 //                   .byteenable
		.avs_readdatavalid ()                                                                                 //        (terminated)
	);

	hls_sim_mm_agent_dpi_bfm #(
		.AV_ADDRESS_W               (64),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (8),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.COMPONENT_NAME             ("relu2"),
		.INTERFACE_ID               (0)
	) mm_agent_dpi_bfm_relu2_avmm_0_rw_inst (
		.do_bind           (relu2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),   //   dpi_control_bind.conduit
		.enable            (relu2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // dpi_control_enable.conduit
		.clock             (clock_reset_inst_clock_clk),                                                      //              clock.clk
		.reset_n           (clock_reset_inst_reset_reset),                                                    //              reset.reset_n
		.avs_writedata     (relu2_inst_avmm_0_rw_writedata),                                                  //                 s0.writedata
		.avs_readdata      (relu2_inst_avmm_0_rw_readdata),                                                   //                   .readdata
		.avs_address       (relu2_inst_avmm_0_rw_address),                                                    //                   .address
		.avs_write         (relu2_inst_avmm_0_rw_write),                                                      //                   .write
		.avs_read          (relu2_inst_avmm_0_rw_read),                                                       //                   .read
		.avs_byteenable    (relu2_inst_avmm_0_rw_byteenable),                                                 //                   .byteenable
		.avs_readdatavalid ()                                                                                 //        (terminated)
	);

	hls_sim_mm_agent_dpi_bfm #(
		.AV_ADDRESS_W               (64),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (8),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.COMPONENT_NAME             ("relu3"),
		.INTERFACE_ID               (0)
	) mm_agent_dpi_bfm_relu3_avmm_0_rw_inst (
		.do_bind           (relu3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),   //   dpi_control_bind.conduit
		.enable            (relu3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // dpi_control_enable.conduit
		.clock             (clock_reset_inst_clock_clk),                                                      //              clock.clk
		.reset_n           (clock_reset_inst_reset_reset),                                                    //              reset.reset_n
		.avs_writedata     (relu3_inst_avmm_0_rw_writedata),                                                  //                 s0.writedata
		.avs_readdata      (relu3_inst_avmm_0_rw_readdata),                                                   //                   .readdata
		.avs_address       (relu3_inst_avmm_0_rw_address),                                                    //                   .address
		.avs_write         (relu3_inst_avmm_0_rw_write),                                                      //                   .write
		.avs_read          (relu3_inst_avmm_0_rw_read),                                                       //                   .read
		.avs_byteenable    (relu3_inst_avmm_0_rw_byteenable),                                                 //                   .byteenable
		.avs_readdatavalid ()                                                                                 //        (terminated)
	);

	hls_sim_mm_agent_dpi_bfm #(
		.AV_ADDRESS_W               (64),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (8),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.COMPONENT_NAME             ("relu4"),
		.INTERFACE_ID               (0)
	) mm_agent_dpi_bfm_relu4_avmm_0_rw_inst (
		.do_bind           (relu4_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),   //   dpi_control_bind.conduit
		.enable            (relu4_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // dpi_control_enable.conduit
		.clock             (clock_reset_inst_clock_clk),                                                      //              clock.clk
		.reset_n           (clock_reset_inst_reset_reset),                                                    //              reset.reset_n
		.avs_writedata     (relu4_inst_avmm_0_rw_writedata),                                                  //                 s0.writedata
		.avs_readdata      (relu4_inst_avmm_0_rw_readdata),                                                   //                   .readdata
		.avs_address       (relu4_inst_avmm_0_rw_address),                                                    //                   .address
		.avs_write         (relu4_inst_avmm_0_rw_write),                                                      //                   .write
		.avs_read          (relu4_inst_avmm_0_rw_read),                                                       //                   .read
		.avs_byteenable    (relu4_inst_avmm_0_rw_byteenable),                                                 //                   .byteenable
		.avs_readdatavalid ()                                                                                 //        (terminated)
	);

	hls_sim_mm_agent_dpi_bfm #(
		.AV_ADDRESS_W               (64),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (8),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.COMPONENT_NAME             ("softmax"),
		.INTERFACE_ID               (0)
	) mm_agent_dpi_bfm_softmax_avmm_0_rw_inst (
		.do_bind           (softmax_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),   //   dpi_control_bind.conduit
		.enable            (softmax_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // dpi_control_enable.conduit
		.clock             (clock_reset_inst_clock_clk),                                                        //              clock.clk
		.reset_n           (clock_reset_inst_reset_reset),                                                      //              reset.reset_n
		.avs_writedata     (softmax_inst_avmm_0_rw_writedata),                                                  //                 s0.writedata
		.avs_readdata      (softmax_inst_avmm_0_rw_readdata),                                                   //                   .readdata
		.avs_address       (softmax_inst_avmm_0_rw_address),                                                    //                   .address
		.avs_write         (softmax_inst_avmm_0_rw_write),                                                      //                   .write
		.avs_read          (softmax_inst_avmm_0_rw_read),                                                       //                   .read
		.avs_byteenable    (softmax_inst_avmm_0_rw_byteenable),                                                 //                   .byteenable
		.avs_readdatavalid ()                                                                                   //        (terminated)
	);

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst relu1_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_relu1_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (relu1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (relu1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (relu1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst relu1_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_relu1_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (relu1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (relu1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (relu1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst relu1_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_relu1_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (relu1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (relu1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit)  // out_conduit_1.conduit
	);

	tb_relu1_inst relu1_inst (
		.avmm_0_rw_address    (relu1_inst_avmm_0_rw_address),                               // avmm_0_rw.address
		.avmm_0_rw_byteenable (relu1_inst_avmm_0_rw_byteenable),                            //          .byteenable
		.avmm_0_rw_read       (relu1_inst_avmm_0_rw_read),                                  //          .read
		.avmm_0_rw_readdata   (relu1_inst_avmm_0_rw_readdata),                              //          .readdata
		.avmm_0_rw_write      (relu1_inst_avmm_0_rw_write),                                 //          .write
		.avmm_0_rw_writedata  (relu1_inst_avmm_0_rw_writedata),                             //          .writedata
		.start                (component_dpi_controller_relu1_inst_component_call_valid),   //      call.valid
		.busy                 (relu1_inst_call_stall),                                      //          .stall
		.clock                (clock_reset_inst_clock_clk),                                 //     clock.clk
		.in0                  (stream_source_dpi_bfm_relu1_in0_inst_source_data_data),      //       in0.data
		.out0                 (stream_source_dpi_bfm_relu1_out0_inst_source_data_data),     //      out0.data
		.resetn               (clock_reset_inst_reset_reset),                               //     reset.reset_n
		.done                 (relu1_inst_return_valid),                                    //    return.valid
		.stall                (component_dpi_controller_relu1_inst_component_return_stall)  //          .stall
	);

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst relu2_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_relu2_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (relu2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (relu2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (relu2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst relu2_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_relu2_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (relu2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (relu2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (relu2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst relu2_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_relu2_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (relu2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (relu2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit)  // out_conduit_1.conduit
	);

	tb_relu2_inst relu2_inst (
		.avmm_0_rw_address    (relu2_inst_avmm_0_rw_address),                               // avmm_0_rw.address
		.avmm_0_rw_byteenable (relu2_inst_avmm_0_rw_byteenable),                            //          .byteenable
		.avmm_0_rw_read       (relu2_inst_avmm_0_rw_read),                                  //          .read
		.avmm_0_rw_readdata   (relu2_inst_avmm_0_rw_readdata),                              //          .readdata
		.avmm_0_rw_write      (relu2_inst_avmm_0_rw_write),                                 //          .write
		.avmm_0_rw_writedata  (relu2_inst_avmm_0_rw_writedata),                             //          .writedata
		.start                (component_dpi_controller_relu2_inst_component_call_valid),   //      call.valid
		.busy                 (relu2_inst_call_stall),                                      //          .stall
		.clock                (clock_reset_inst_clock_clk),                                 //     clock.clk
		.in0                  (stream_source_dpi_bfm_relu2_in0_inst_source_data_data),      //       in0.data
		.out0                 (stream_source_dpi_bfm_relu2_out0_inst_source_data_data),     //      out0.data
		.resetn               (clock_reset_inst_reset_reset),                               //     reset.reset_n
		.done                 (relu2_inst_return_valid),                                    //    return.valid
		.stall                (component_dpi_controller_relu2_inst_component_return_stall)  //          .stall
	);

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst relu3_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_relu3_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (relu3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (relu3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (relu3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst relu3_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_relu3_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (relu3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (relu3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (relu3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst relu3_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_relu3_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (relu3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (relu3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit)  // out_conduit_1.conduit
	);

	tb_relu3_inst relu3_inst (
		.avmm_0_rw_address    (relu3_inst_avmm_0_rw_address),                               // avmm_0_rw.address
		.avmm_0_rw_byteenable (relu3_inst_avmm_0_rw_byteenable),                            //          .byteenable
		.avmm_0_rw_read       (relu3_inst_avmm_0_rw_read),                                  //          .read
		.avmm_0_rw_readdata   (relu3_inst_avmm_0_rw_readdata),                              //          .readdata
		.avmm_0_rw_write      (relu3_inst_avmm_0_rw_write),                                 //          .write
		.avmm_0_rw_writedata  (relu3_inst_avmm_0_rw_writedata),                             //          .writedata
		.start                (component_dpi_controller_relu3_inst_component_call_valid),   //      call.valid
		.busy                 (relu3_inst_call_stall),                                      //          .stall
		.clock                (clock_reset_inst_clock_clk),                                 //     clock.clk
		.in0                  (stream_source_dpi_bfm_relu3_in0_inst_source_data_data),      //       in0.data
		.out0                 (stream_source_dpi_bfm_relu3_out0_inst_source_data_data),     //      out0.data
		.resetn               (clock_reset_inst_reset_reset),                               //     reset.reset_n
		.done                 (relu3_inst_return_valid),                                    //    return.valid
		.stall                (component_dpi_controller_relu3_inst_component_return_stall)  //          .stall
	);

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst relu4_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_relu4_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (relu4_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (relu4_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (relu4_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst relu4_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_relu4_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (relu4_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (relu4_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (relu4_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst relu4_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_relu4_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (relu4_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (relu4_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit)  // out_conduit_1.conduit
	);

	tb_relu4_inst relu4_inst (
		.avmm_0_rw_address    (relu4_inst_avmm_0_rw_address),                               // avmm_0_rw.address
		.avmm_0_rw_byteenable (relu4_inst_avmm_0_rw_byteenable),                            //          .byteenable
		.avmm_0_rw_read       (relu4_inst_avmm_0_rw_read),                                  //          .read
		.avmm_0_rw_readdata   (relu4_inst_avmm_0_rw_readdata),                              //          .readdata
		.avmm_0_rw_write      (relu4_inst_avmm_0_rw_write),                                 //          .write
		.avmm_0_rw_writedata  (relu4_inst_avmm_0_rw_writedata),                             //          .writedata
		.start                (component_dpi_controller_relu4_inst_component_call_valid),   //      call.valid
		.busy                 (relu4_inst_call_stall),                                      //          .stall
		.clock                (clock_reset_inst_clock_clk),                                 //     clock.clk
		.in0                  (stream_source_dpi_bfm_relu4_in0_inst_source_data_data),      //       in0.data
		.out0                 (stream_source_dpi_bfm_relu4_out0_inst_source_data_data),     //      out0.data
		.resetn               (clock_reset_inst_reset_reset),                               //     reset.reset_n
		.done                 (relu4_inst_return_valid),                                    //    return.valid
		.stall                (component_dpi_controller_relu4_inst_component_return_stall)  //          .stall
	);

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst softmax_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_softmax_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (softmax_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (softmax_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (softmax_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_bind_conduit_fanout_inst softmax_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_softmax_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (softmax_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (softmax_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (softmax_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst softmax_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_softmax_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (softmax_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (softmax_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit)  // out_conduit_1.conduit
	);

	tb_softmax_inst softmax_inst (
		.avmm_0_rw_address    (softmax_inst_avmm_0_rw_address),                               // avmm_0_rw.address
		.avmm_0_rw_byteenable (softmax_inst_avmm_0_rw_byteenable),                            //          .byteenable
		.avmm_0_rw_read       (softmax_inst_avmm_0_rw_read),                                  //          .read
		.avmm_0_rw_readdata   (softmax_inst_avmm_0_rw_readdata),                              //          .readdata
		.avmm_0_rw_write      (softmax_inst_avmm_0_rw_write),                                 //          .write
		.avmm_0_rw_writedata  (softmax_inst_avmm_0_rw_writedata),                             //          .writedata
		.start                (component_dpi_controller_softmax_inst_component_call_valid),   //      call.valid
		.busy                 (softmax_inst_call_stall),                                      //          .stall
		.clock                (clock_reset_inst_clock_clk),                                   //     clock.clk
		.in0                  (stream_source_dpi_bfm_softmax_in0_inst_source_data_data),      //       in0.data
		.out0                 (stream_source_dpi_bfm_softmax_out0_inst_source_data_data),     //      out0.data
		.resetn               (clock_reset_inst_reset_reset),                                 //     reset.reset_n
		.done                 (softmax_inst_return_valid),                                    //    return.valid
		.stall                (component_dpi_controller_softmax_inst_component_return_stall)  //          .stall
	);

	tb_split_component_start_inst split_component_start_inst (
		.in_conduit     (main_dpi_controller_inst_component_enabled_conduit), //     in_conduit.conduit
		.out_conduit_0  (split_component_start_inst_out_conduit_0_conduit),   //  out_conduit_0.conduit
		.out_conduit_1  (split_component_start_inst_out_conduit_1_conduit),   //  out_conduit_1.conduit
		.out_conduit_2  (split_component_start_inst_out_conduit_2_conduit),   //  out_conduit_2.conduit
		.out_conduit_3  (split_component_start_inst_out_conduit_3_conduit),   //  out_conduit_3.conduit
		.out_conduit_4  (split_component_start_inst_out_conduit_4_conduit),   //  out_conduit_4.conduit
		.out_conduit_5  (split_component_start_inst_out_conduit_5_conduit),   //  out_conduit_5.conduit
		.out_conduit_6  (split_component_start_inst_out_conduit_6_conduit),   //  out_conduit_6.conduit
		.out_conduit_7  (split_component_start_inst_out_conduit_7_conduit),   //  out_conduit_7.conduit
		.out_conduit_8  (split_component_start_inst_out_conduit_8_conduit),   //  out_conduit_8.conduit
		.out_conduit_9  (split_component_start_inst_out_conduit_9_conduit),   //  out_conduit_9.conduit
		.out_conduit_10 (split_component_start_inst_out_conduit_10_conduit)   // out_conduit_10.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("avgpooling1"),
		.INTERFACE_NAME                  ("in"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_avgpooling1_in0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                    //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                  //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                  //            clock2x.clk
		.do_bind      (avgpooling1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //   dpi_control_bind.conduit
		.enable       (avgpooling1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_avgpooling1_in0_inst_source_data_data),                                   //        source_data.data
		.source_ready (avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                               //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("avgpooling1"),
		.INTERFACE_NAME                  ("out"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_avgpooling1_out0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                    //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                  //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                  //            clock2x.clk
		.do_bind      (avgpooling1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //   dpi_control_bind.conduit
		.enable       (avgpooling1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_avgpooling1_out0_inst_source_data_data),                                  //        source_data.data
		.source_ready (avgpooling1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //       source_ready.conduit
		.source_valid ()                                                                                               //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("avgpooling2"),
		.INTERFACE_NAME                  ("in"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_avgpooling2_in0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                    //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                  //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                  //            clock2x.clk
		.do_bind      (avgpooling2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //   dpi_control_bind.conduit
		.enable       (avgpooling2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_avgpooling2_in0_inst_source_data_data),                                   //        source_data.data
		.source_ready (avgpooling2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                               //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("avgpooling2"),
		.INTERFACE_NAME                  ("out"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_avgpooling2_out0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                    //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                  //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                  //            clock2x.clk
		.do_bind      (avgpooling2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //   dpi_control_bind.conduit
		.enable       (avgpooling2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_avgpooling2_out0_inst_source_data_data),                                  //        source_data.data
		.source_ready (avgpooling2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //       source_ready.conduit
		.source_valid ()                                                                                               //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("conv1"),
		.INTERFACE_NAME                  ("bias"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_conv1_bias_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //   dpi_control_bind.conduit
		.enable       (conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_conv1_bias_inst_source_data_data),                                  //        source_data.data
		.source_ready (conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("conv1"),
		.INTERFACE_NAME                  ("in"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_conv1_in0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //   dpi_control_bind.conduit
		.enable       (conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_conv1_in0_inst_source_data_data),                                   //        source_data.data
		.source_ready (conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("conv1"),
		.INTERFACE_NAME                  ("kernel"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_conv1_kernel_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit),           //   dpi_control_bind.conduit
		.enable       (conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_conv1_kernel_inst_source_data_data),                                //        source_data.data
		.source_ready (conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("conv1"),
		.INTERFACE_NAME                  ("out"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_conv1_out0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (conv1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit),           //   dpi_control_bind.conduit
		.enable       (conv1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_conv1_out0_inst_source_data_data),                                  //        source_data.data
		.source_ready (conv1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("conv2"),
		.INTERFACE_NAME                  ("bias"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_conv2_bias_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //   dpi_control_bind.conduit
		.enable       (conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_conv2_bias_inst_source_data_data),                                  //        source_data.data
		.source_ready (conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("conv2"),
		.INTERFACE_NAME                  ("in"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_conv2_in0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //   dpi_control_bind.conduit
		.enable       (conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_conv2_in0_inst_source_data_data),                                   //        source_data.data
		.source_ready (conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("conv2"),
		.INTERFACE_NAME                  ("kernel"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_conv2_kernel_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit),           //   dpi_control_bind.conduit
		.enable       (conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_conv2_kernel_inst_source_data_data),                                //        source_data.data
		.source_ready (conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("conv2"),
		.INTERFACE_NAME                  ("out"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_conv2_out0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (conv2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit),           //   dpi_control_bind.conduit
		.enable       (conv2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_conv2_out0_inst_source_data_data),                                  //        source_data.data
		.source_ready (conv2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("fc1"),
		.INTERFACE_NAME                  ("bias"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_fc1_bias_inst (
		.clock        (clock_reset_inst_clock_clk),                                                            //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                          //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                          //            clock2x.clk
		.do_bind      (fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //   dpi_control_bind.conduit
		.enable       (fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_fc1_bias_inst_source_data_data),                                  //        source_data.data
		.source_ready (fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                       //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("fc1"),
		.INTERFACE_NAME                  ("in"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_fc1_in0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                            //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                          //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                          //            clock2x.clk
		.do_bind      (fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //   dpi_control_bind.conduit
		.enable       (fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_fc1_in0_inst_source_data_data),                                   //        source_data.data
		.source_ready (fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //       source_ready.conduit
		.source_valid ()                                                                                       //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("fc1"),
		.INTERFACE_NAME                  ("out"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_fc1_out0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                            //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                          //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                          //            clock2x.clk
		.do_bind      (fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit),           //   dpi_control_bind.conduit
		.enable       (fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_fc1_out0_inst_source_data_data),                                  //        source_data.data
		.source_ready (fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit), //       source_ready.conduit
		.source_valid ()                                                                                       //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("fc1"),
		.INTERFACE_NAME                  ("weights"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_fc1_weights_inst (
		.clock        (clock_reset_inst_clock_clk),                                                            //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                          //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                          //            clock2x.clk
		.do_bind      (fc1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit),           //   dpi_control_bind.conduit
		.enable       (fc1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_fc1_weights_inst_source_data_data),                               //        source_data.data
		.source_ready (fc1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit), //       source_ready.conduit
		.source_valid ()                                                                                       //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("fc3"),
		.INTERFACE_NAME                  ("bias"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_fc3_bias_inst (
		.clock        (clock_reset_inst_clock_clk),                                                            //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                          //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                          //            clock2x.clk
		.do_bind      (fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //   dpi_control_bind.conduit
		.enable       (fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_fc3_bias_inst_source_data_data),                                  //        source_data.data
		.source_ready (fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                       //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("fc3"),
		.INTERFACE_NAME                  ("in"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_fc3_in0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                            //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                          //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                          //            clock2x.clk
		.do_bind      (fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //   dpi_control_bind.conduit
		.enable       (fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_fc3_in0_inst_source_data_data),                                   //        source_data.data
		.source_ready (fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //       source_ready.conduit
		.source_valid ()                                                                                       //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("fc3"),
		.INTERFACE_NAME                  ("out"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_fc3_out0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                            //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                          //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                          //            clock2x.clk
		.do_bind      (fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit),           //   dpi_control_bind.conduit
		.enable       (fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_fc3_out0_inst_source_data_data),                                  //        source_data.data
		.source_ready (fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit), //       source_ready.conduit
		.source_valid ()                                                                                       //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("fc3"),
		.INTERFACE_NAME                  ("weights"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_fc3_weights_inst (
		.clock        (clock_reset_inst_clock_clk),                                                            //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                          //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                          //            clock2x.clk
		.do_bind      (fc3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit),           //   dpi_control_bind.conduit
		.enable       (fc3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_fc3_weights_inst_source_data_data),                               //        source_data.data
		.source_ready (fc3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit), //       source_ready.conduit
		.source_valid ()                                                                                       //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("relu1"),
		.INTERFACE_NAME                  ("in"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_relu1_in0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (relu1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //   dpi_control_bind.conduit
		.enable       (relu1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_relu1_in0_inst_source_data_data),                                   //        source_data.data
		.source_ready (relu1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("relu1"),
		.INTERFACE_NAME                  ("out"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_relu1_out0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (relu1_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //   dpi_control_bind.conduit
		.enable       (relu1_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_relu1_out0_inst_source_data_data),                                  //        source_data.data
		.source_ready (relu1_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("relu2"),
		.INTERFACE_NAME                  ("in"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_relu2_in0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (relu2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //   dpi_control_bind.conduit
		.enable       (relu2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_relu2_in0_inst_source_data_data),                                   //        source_data.data
		.source_ready (relu2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("relu2"),
		.INTERFACE_NAME                  ("out"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_relu2_out0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (relu2_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //   dpi_control_bind.conduit
		.enable       (relu2_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_relu2_out0_inst_source_data_data),                                  //        source_data.data
		.source_ready (relu2_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("relu3"),
		.INTERFACE_NAME                  ("in"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_relu3_in0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (relu3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //   dpi_control_bind.conduit
		.enable       (relu3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_relu3_in0_inst_source_data_data),                                   //        source_data.data
		.source_ready (relu3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("relu3"),
		.INTERFACE_NAME                  ("out"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_relu3_out0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (relu3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //   dpi_control_bind.conduit
		.enable       (relu3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_relu3_out0_inst_source_data_data),                                  //        source_data.data
		.source_ready (relu3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("relu4"),
		.INTERFACE_NAME                  ("in"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_relu4_in0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (relu4_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //   dpi_control_bind.conduit
		.enable       (relu4_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_relu4_in0_inst_source_data_data),                                   //        source_data.data
		.source_ready (relu4_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("relu4"),
		.INTERFACE_NAME                  ("out"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_relu4_out0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                              //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                            //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                            //            clock2x.clk
		.do_bind      (relu4_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //   dpi_control_bind.conduit
		.enable       (relu4_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_relu4_out0_inst_source_data_data),                                  //        source_data.data
		.source_ready (relu4_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //       source_ready.conduit
		.source_valid ()                                                                                         //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("softmax"),
		.INTERFACE_NAME                  ("in"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_softmax_in0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                              //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                              //            clock2x.clk
		.do_bind      (softmax_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //   dpi_control_bind.conduit
		.enable       (softmax_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_softmax_in0_inst_source_data_data),                                   //        source_data.data
		.source_ready (softmax_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                           //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("softmax"),
		.INTERFACE_NAME                  ("out"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_softmax_out0_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                              //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                              //            clock2x.clk
		.do_bind      (softmax_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //   dpi_control_bind.conduit
		.enable       (softmax_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_softmax_out0_inst_source_data_data),                                  //        source_data.data
		.source_ready (softmax_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //       source_ready.conduit
		.source_valid ()                                                                                           //             source.conduit
	);

	tb_irq_mapper irq_mapper (
		.clk        (clock_reset_inst_clock_clk),                                  //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                               // clk_reset.reset
		.sender_irq (component_dpi_controller_avgpooling1_inst_component_irq_irq)  //    sender.irq
	);

	tb_irq_mapper irq_mapper_001 (
		.clk        (clock_reset_inst_clock_clk),                                  //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                               // clk_reset.reset
		.sender_irq (component_dpi_controller_avgpooling2_inst_component_irq_irq)  //    sender.irq
	);

	tb_irq_mapper irq_mapper_002 (
		.clk        (clock_reset_inst_clock_clk),                            //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                         // clk_reset.reset
		.sender_irq (component_dpi_controller_conv1_inst_component_irq_irq)  //    sender.irq
	);

	tb_irq_mapper irq_mapper_003 (
		.clk        (clock_reset_inst_clock_clk),                            //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                         // clk_reset.reset
		.sender_irq (component_dpi_controller_conv2_inst_component_irq_irq)  //    sender.irq
	);

	tb_irq_mapper irq_mapper_004 (
		.clk        (clock_reset_inst_clock_clk),                          //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                       // clk_reset.reset
		.sender_irq (component_dpi_controller_fc1_inst_component_irq_irq)  //    sender.irq
	);

	tb_irq_mapper irq_mapper_005 (
		.clk        (clock_reset_inst_clock_clk),                          //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                       // clk_reset.reset
		.sender_irq (component_dpi_controller_fc3_inst_component_irq_irq)  //    sender.irq
	);

	tb_irq_mapper irq_mapper_006 (
		.clk        (clock_reset_inst_clock_clk),                            //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                         // clk_reset.reset
		.sender_irq (component_dpi_controller_relu1_inst_component_irq_irq)  //    sender.irq
	);

	tb_irq_mapper irq_mapper_007 (
		.clk        (clock_reset_inst_clock_clk),                            //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                         // clk_reset.reset
		.sender_irq (component_dpi_controller_relu2_inst_component_irq_irq)  //    sender.irq
	);

	tb_irq_mapper irq_mapper_008 (
		.clk        (clock_reset_inst_clock_clk),                            //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                         // clk_reset.reset
		.sender_irq (component_dpi_controller_relu3_inst_component_irq_irq)  //    sender.irq
	);

	tb_irq_mapper irq_mapper_009 (
		.clk        (clock_reset_inst_clock_clk),                            //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                         // clk_reset.reset
		.sender_irq (component_dpi_controller_relu4_inst_component_irq_irq)  //    sender.irq
	);

	tb_irq_mapper irq_mapper_010 (
		.clk        (clock_reset_inst_clock_clk),                              //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                           // clk_reset.reset
		.sender_irq (component_dpi_controller_softmax_inst_component_irq_irq)  //    sender.irq
	);

endmodule
